magic
tech gf180mcuC
magscale 1 10
timestamp 1670279682
<< metal1 >>
rect 35970 57038 35982 57090
rect 36034 57087 36046 57090
rect 37090 57087 37102 57090
rect 36034 57041 37102 57087
rect 36034 57038 36046 57041
rect 37090 57038 37102 57041
rect 37154 57038 37166 57090
rect 53890 56926 53902 56978
rect 53954 56975 53966 56978
rect 54674 56975 54686 56978
rect 53954 56929 54686 56975
rect 53954 56926 53966 56929
rect 54674 56926 54686 56929
rect 54738 56926 54750 56978
rect 44482 56814 44494 56866
rect 44546 56863 44558 56866
rect 45602 56863 45614 56866
rect 44546 56817 45614 56863
rect 44546 56814 44558 56817
rect 45602 56814 45614 56817
rect 45666 56814 45678 56866
rect 34626 56702 34638 56754
rect 34690 56751 34702 56754
rect 35186 56751 35198 56754
rect 34690 56705 35198 56751
rect 34690 56702 34702 56705
rect 35186 56702 35198 56705
rect 35250 56702 35262 56754
rect 44034 56702 44046 56754
rect 44098 56751 44110 56754
rect 44930 56751 44942 56754
rect 44098 56705 44942 56751
rect 44098 56702 44110 56705
rect 44930 56702 44942 56705
rect 44994 56702 45006 56754
rect 45826 56702 45838 56754
rect 45890 56751 45902 56754
rect 46946 56751 46958 56754
rect 45890 56705 46958 56751
rect 45890 56702 45902 56705
rect 46946 56702 46958 56705
rect 47010 56702 47022 56754
rect 48738 56702 48750 56754
rect 48802 56751 48814 56754
rect 49522 56751 49534 56754
rect 48802 56705 49534 56751
rect 48802 56702 48814 56705
rect 49522 56702 49534 56705
rect 49586 56702 49598 56754
rect 49858 56702 49870 56754
rect 49922 56751 49934 56754
rect 50866 56751 50878 56754
rect 49922 56705 50878 56751
rect 49922 56702 49934 56705
rect 50866 56702 50878 56705
rect 50930 56702 50942 56754
rect 52546 56702 52558 56754
rect 52610 56751 52622 56754
rect 53330 56751 53342 56754
rect 52610 56705 53342 56751
rect 52610 56702 52622 56705
rect 53330 56702 53342 56705
rect 53394 56702 53406 56754
rect 20626 56590 20638 56642
rect 20690 56639 20702 56642
rect 21186 56639 21198 56642
rect 20690 56593 21198 56639
rect 20690 56590 20702 56593
rect 21186 56590 21198 56593
rect 21250 56590 21262 56642
rect 32386 56590 32398 56642
rect 32450 56639 32462 56642
rect 33170 56639 33182 56642
rect 32450 56593 33182 56639
rect 32450 56590 32462 56593
rect 33170 56590 33182 56593
rect 33234 56590 33246 56642
rect 33730 56590 33742 56642
rect 33794 56639 33806 56642
rect 34514 56639 34526 56642
rect 33794 56593 34526 56639
rect 33794 56590 33806 56593
rect 34514 56590 34526 56593
rect 34578 56590 34590 56642
rect 37874 56590 37886 56642
rect 37938 56639 37950 56642
rect 38434 56639 38446 56642
rect 37938 56593 38446 56639
rect 37938 56590 37950 56593
rect 38434 56590 38446 56593
rect 38498 56590 38510 56642
rect 39218 56590 39230 56642
rect 39282 56639 39294 56642
rect 39778 56639 39790 56642
rect 39282 56593 39790 56639
rect 39282 56590 39294 56593
rect 39778 56590 39790 56593
rect 39842 56590 39854 56642
rect 40450 56590 40462 56642
rect 40514 56639 40526 56642
rect 41682 56639 41694 56642
rect 40514 56593 41694 56639
rect 40514 56590 40526 56593
rect 41682 56590 41694 56593
rect 41746 56590 41758 56642
rect 45378 56590 45390 56642
rect 45442 56639 45454 56642
rect 46274 56639 46286 56642
rect 45442 56593 46286 56639
rect 45442 56590 45454 56593
rect 46274 56590 46286 56593
rect 46338 56590 46350 56642
rect 49410 56590 49422 56642
rect 49474 56639 49486 56642
rect 50194 56639 50206 56642
rect 49474 56593 50206 56639
rect 49474 56590 49486 56593
rect 50194 56590 50206 56593
rect 50258 56590 50270 56642
rect 50754 56590 50766 56642
rect 50818 56639 50830 56642
rect 51538 56639 51550 56642
rect 50818 56593 51550 56639
rect 50818 56590 50830 56593
rect 51538 56590 51550 56593
rect 51602 56590 51614 56642
rect 52098 56590 52110 56642
rect 52162 56639 52174 56642
rect 52770 56639 52782 56642
rect 52162 56593 52782 56639
rect 52162 56590 52174 56593
rect 52770 56590 52782 56593
rect 52834 56590 52846 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 4958 56306 5010 56318
rect 4958 56242 5010 56254
rect 6190 56306 6242 56318
rect 6190 56242 6242 56254
rect 6862 56306 6914 56318
rect 6862 56242 6914 56254
rect 7534 56306 7586 56318
rect 7534 56242 7586 56254
rect 8206 56306 8258 56318
rect 8206 56242 8258 56254
rect 8878 56306 8930 56318
rect 8878 56242 8930 56254
rect 10110 56306 10162 56318
rect 10110 56242 10162 56254
rect 10782 56306 10834 56318
rect 10782 56242 10834 56254
rect 12126 56306 12178 56318
rect 12126 56242 12178 56254
rect 14702 56306 14754 56318
rect 14702 56242 14754 56254
rect 16046 56306 16098 56318
rect 16046 56242 16098 56254
rect 17838 56306 17890 56318
rect 17838 56242 17890 56254
rect 19182 56306 19234 56318
rect 19182 56242 19234 56254
rect 19966 56306 20018 56318
rect 19966 56242 20018 56254
rect 21758 56306 21810 56318
rect 21758 56242 21810 56254
rect 23102 56306 23154 56318
rect 23102 56242 23154 56254
rect 24446 56306 24498 56318
rect 24446 56242 24498 56254
rect 25678 56306 25730 56318
rect 25678 56242 25730 56254
rect 27022 56306 27074 56318
rect 27022 56242 27074 56254
rect 28366 56306 28418 56318
rect 28366 56242 28418 56254
rect 29934 56306 29986 56318
rect 29934 56242 29986 56254
rect 31278 56306 31330 56318
rect 31278 56242 31330 56254
rect 33182 56306 33234 56318
rect 33182 56242 33234 56254
rect 34526 56306 34578 56318
rect 34526 56242 34578 56254
rect 35198 56306 35250 56318
rect 35198 56242 35250 56254
rect 37102 56306 37154 56318
rect 37102 56242 37154 56254
rect 37774 56306 37826 56318
rect 37774 56242 37826 56254
rect 38446 56306 38498 56318
rect 38446 56242 38498 56254
rect 39118 56306 39170 56318
rect 39118 56242 39170 56254
rect 39790 56306 39842 56318
rect 39790 56242 39842 56254
rect 41022 56306 41074 56318
rect 41022 56242 41074 56254
rect 41694 56306 41746 56318
rect 41694 56242 41746 56254
rect 42366 56306 42418 56318
rect 42366 56242 42418 56254
rect 43038 56306 43090 56318
rect 43038 56242 43090 56254
rect 43710 56306 43762 56318
rect 43710 56242 43762 56254
rect 44942 56306 44994 56318
rect 44942 56242 44994 56254
rect 45614 56306 45666 56318
rect 45614 56242 45666 56254
rect 46286 56306 46338 56318
rect 46286 56242 46338 56254
rect 46958 56306 47010 56318
rect 46958 56242 47010 56254
rect 48862 56306 48914 56318
rect 48862 56242 48914 56254
rect 49534 56306 49586 56318
rect 49534 56242 49586 56254
rect 50206 56306 50258 56318
rect 50206 56242 50258 56254
rect 50878 56306 50930 56318
rect 50878 56242 50930 56254
rect 51550 56306 51602 56318
rect 51550 56242 51602 56254
rect 52782 56306 52834 56318
rect 52782 56242 52834 56254
rect 53454 56306 53506 56318
rect 53454 56242 53506 56254
rect 54126 56306 54178 56318
rect 54126 56242 54178 56254
rect 55470 56306 55522 56318
rect 55470 56242 55522 56254
rect 11454 56194 11506 56206
rect 11454 56130 11506 56142
rect 35870 56194 35922 56206
rect 35870 56130 35922 56142
rect 47630 56194 47682 56206
rect 47630 56130 47682 56142
rect 54798 56194 54850 56206
rect 54798 56130 54850 56142
rect 12798 55970 12850 55982
rect 12798 55906 12850 55918
rect 14030 55970 14082 55982
rect 14030 55906 14082 55918
rect 15374 55970 15426 55982
rect 15374 55906 15426 55918
rect 16718 55970 16770 55982
rect 16718 55906 16770 55918
rect 18510 55970 18562 55982
rect 18510 55906 18562 55918
rect 20638 55970 20690 55982
rect 20638 55906 20690 55918
rect 22542 55970 22594 55982
rect 22542 55906 22594 55918
rect 23886 55970 23938 55982
rect 23886 55906 23938 55918
rect 26462 55970 26514 55982
rect 26462 55906 26514 55918
rect 27806 55970 27858 55982
rect 27806 55906 27858 55918
rect 29262 55970 29314 55982
rect 29262 55906 29314 55918
rect 30606 55970 30658 55982
rect 30606 55906 30658 55918
rect 32174 55970 32226 55982
rect 32174 55906 32226 55918
rect 33854 55970 33906 55982
rect 33854 55906 33906 55918
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 20078 55522 20130 55534
rect 20078 55458 20130 55470
rect 25454 55522 25506 55534
rect 25454 55458 25506 55470
rect 5742 55186 5794 55198
rect 5742 55122 5794 55134
rect 9774 55186 9826 55198
rect 9774 55122 9826 55134
rect 13806 55186 13858 55198
rect 13806 55122 13858 55134
rect 36654 55186 36706 55198
rect 36654 55122 36706 55134
rect 43374 55186 43426 55198
rect 43374 55122 43426 55134
rect 47406 55186 47458 55198
rect 47406 55122 47458 55134
rect 51438 55186 51490 55198
rect 51438 55122 51490 55134
rect 55470 55186 55522 55198
rect 55470 55122 55522 55134
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 35982 57038 36034 57090
rect 37102 57038 37154 57090
rect 53902 56926 53954 56978
rect 54686 56926 54738 56978
rect 44494 56814 44546 56866
rect 45614 56814 45666 56866
rect 34638 56702 34690 56754
rect 35198 56702 35250 56754
rect 44046 56702 44098 56754
rect 44942 56702 44994 56754
rect 45838 56702 45890 56754
rect 46958 56702 47010 56754
rect 48750 56702 48802 56754
rect 49534 56702 49586 56754
rect 49870 56702 49922 56754
rect 50878 56702 50930 56754
rect 52558 56702 52610 56754
rect 53342 56702 53394 56754
rect 20638 56590 20690 56642
rect 21198 56590 21250 56642
rect 32398 56590 32450 56642
rect 33182 56590 33234 56642
rect 33742 56590 33794 56642
rect 34526 56590 34578 56642
rect 37886 56590 37938 56642
rect 38446 56590 38498 56642
rect 39230 56590 39282 56642
rect 39790 56590 39842 56642
rect 40462 56590 40514 56642
rect 41694 56590 41746 56642
rect 45390 56590 45442 56642
rect 46286 56590 46338 56642
rect 49422 56590 49474 56642
rect 50206 56590 50258 56642
rect 50766 56590 50818 56642
rect 51550 56590 51602 56642
rect 52110 56590 52162 56642
rect 52782 56590 52834 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 4958 56254 5010 56306
rect 6190 56254 6242 56306
rect 6862 56254 6914 56306
rect 7534 56254 7586 56306
rect 8206 56254 8258 56306
rect 8878 56254 8930 56306
rect 10110 56254 10162 56306
rect 10782 56254 10834 56306
rect 12126 56254 12178 56306
rect 14702 56254 14754 56306
rect 16046 56254 16098 56306
rect 17838 56254 17890 56306
rect 19182 56254 19234 56306
rect 19966 56254 20018 56306
rect 21758 56254 21810 56306
rect 23102 56254 23154 56306
rect 24446 56254 24498 56306
rect 25678 56254 25730 56306
rect 27022 56254 27074 56306
rect 28366 56254 28418 56306
rect 29934 56254 29986 56306
rect 31278 56254 31330 56306
rect 33182 56254 33234 56306
rect 34526 56254 34578 56306
rect 35198 56254 35250 56306
rect 37102 56254 37154 56306
rect 37774 56254 37826 56306
rect 38446 56254 38498 56306
rect 39118 56254 39170 56306
rect 39790 56254 39842 56306
rect 41022 56254 41074 56306
rect 41694 56254 41746 56306
rect 42366 56254 42418 56306
rect 43038 56254 43090 56306
rect 43710 56254 43762 56306
rect 44942 56254 44994 56306
rect 45614 56254 45666 56306
rect 46286 56254 46338 56306
rect 46958 56254 47010 56306
rect 48862 56254 48914 56306
rect 49534 56254 49586 56306
rect 50206 56254 50258 56306
rect 50878 56254 50930 56306
rect 51550 56254 51602 56306
rect 52782 56254 52834 56306
rect 53454 56254 53506 56306
rect 54126 56254 54178 56306
rect 55470 56254 55522 56306
rect 11454 56142 11506 56194
rect 35870 56142 35922 56194
rect 47630 56142 47682 56194
rect 54798 56142 54850 56194
rect 12798 55918 12850 55970
rect 14030 55918 14082 55970
rect 15374 55918 15426 55970
rect 16718 55918 16770 55970
rect 18510 55918 18562 55970
rect 20638 55918 20690 55970
rect 22542 55918 22594 55970
rect 23886 55918 23938 55970
rect 26462 55918 26514 55970
rect 27806 55918 27858 55970
rect 29262 55918 29314 55970
rect 30606 55918 30658 55970
rect 32174 55918 32226 55970
rect 33854 55918 33906 55970
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 20078 55470 20130 55522
rect 25454 55470 25506 55522
rect 5742 55134 5794 55186
rect 9774 55134 9826 55186
rect 13806 55134 13858 55186
rect 36654 55134 36706 55186
rect 43374 55134 43426 55186
rect 47406 55134 47458 55186
rect 51438 55134 51490 55186
rect 55470 55134 55522 55186
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 4592 59200 4704 60000
rect 5040 59200 5152 60000
rect 5488 59200 5600 60000
rect 5936 59200 6048 60000
rect 6384 59200 6496 60000
rect 6832 59200 6944 60000
rect 7280 59200 7392 60000
rect 7728 59200 7840 60000
rect 8176 59200 8288 60000
rect 8624 59200 8736 60000
rect 9072 59200 9184 60000
rect 9520 59200 9632 60000
rect 9968 59200 10080 60000
rect 10416 59200 10528 60000
rect 10864 59200 10976 60000
rect 11312 59200 11424 60000
rect 11760 59200 11872 60000
rect 12208 59200 12320 60000
rect 12656 59200 12768 60000
rect 13104 59200 13216 60000
rect 13552 59200 13664 60000
rect 14000 59200 14112 60000
rect 14448 59200 14560 60000
rect 14896 59200 15008 60000
rect 15344 59200 15456 60000
rect 15792 59200 15904 60000
rect 16240 59200 16352 60000
rect 16688 59200 16800 60000
rect 17136 59200 17248 60000
rect 17584 59200 17696 60000
rect 18032 59200 18144 60000
rect 18480 59200 18592 60000
rect 18928 59200 19040 60000
rect 19376 59200 19488 60000
rect 19824 59200 19936 60000
rect 20272 59200 20384 60000
rect 20720 59200 20832 60000
rect 21168 59200 21280 60000
rect 21616 59200 21728 60000
rect 22064 59200 22176 60000
rect 22512 59200 22624 60000
rect 22960 59200 23072 60000
rect 23408 59200 23520 60000
rect 23856 59200 23968 60000
rect 24304 59200 24416 60000
rect 24752 59200 24864 60000
rect 25200 59200 25312 60000
rect 25648 59200 25760 60000
rect 26096 59200 26208 60000
rect 26544 59200 26656 60000
rect 26992 59200 27104 60000
rect 27440 59200 27552 60000
rect 27888 59200 28000 60000
rect 28336 59200 28448 60000
rect 28784 59200 28896 60000
rect 29232 59200 29344 60000
rect 29680 59200 29792 60000
rect 30128 59200 30240 60000
rect 30576 59200 30688 60000
rect 31024 59200 31136 60000
rect 31472 59200 31584 60000
rect 31920 59200 32032 60000
rect 32368 59200 32480 60000
rect 32816 59200 32928 60000
rect 33264 59200 33376 60000
rect 33712 59200 33824 60000
rect 34160 59200 34272 60000
rect 34608 59200 34720 60000
rect 35056 59200 35168 60000
rect 35504 59200 35616 60000
rect 35952 59200 36064 60000
rect 36400 59200 36512 60000
rect 36848 59200 36960 60000
rect 37296 59200 37408 60000
rect 37744 59200 37856 60000
rect 38192 59200 38304 60000
rect 38640 59200 38752 60000
rect 39088 59200 39200 60000
rect 39536 59200 39648 60000
rect 39984 59200 40096 60000
rect 40432 59200 40544 60000
rect 40880 59200 40992 60000
rect 41328 59200 41440 60000
rect 41776 59200 41888 60000
rect 42224 59200 42336 60000
rect 42672 59200 42784 60000
rect 43120 59200 43232 60000
rect 43568 59200 43680 60000
rect 44016 59200 44128 60000
rect 44464 59200 44576 60000
rect 44912 59200 45024 60000
rect 45360 59200 45472 60000
rect 45808 59200 45920 60000
rect 46256 59200 46368 60000
rect 46704 59200 46816 60000
rect 47152 59200 47264 60000
rect 47600 59200 47712 60000
rect 48048 59200 48160 60000
rect 48496 59200 48608 60000
rect 48944 59200 49056 60000
rect 49392 59200 49504 60000
rect 49840 59200 49952 60000
rect 50288 59200 50400 60000
rect 50736 59200 50848 60000
rect 51184 59200 51296 60000
rect 51632 59200 51744 60000
rect 52080 59200 52192 60000
rect 52528 59200 52640 60000
rect 52976 59200 53088 60000
rect 53424 59200 53536 60000
rect 53872 59200 53984 60000
rect 54320 59200 54432 60000
rect 54768 59200 54880 60000
rect 55216 59200 55328 60000
rect 4956 56308 5012 56318
rect 5068 56308 5124 59200
rect 4956 56306 5124 56308
rect 4956 56254 4958 56306
rect 5010 56254 5124 56306
rect 4956 56252 5124 56254
rect 4956 56242 5012 56252
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 5516 55188 5572 59200
rect 6188 56308 6244 56318
rect 6412 56308 6468 59200
rect 6188 56306 6468 56308
rect 6188 56254 6190 56306
rect 6242 56254 6468 56306
rect 6188 56252 6468 56254
rect 6860 56306 6916 59200
rect 6860 56254 6862 56306
rect 6914 56254 6916 56306
rect 6188 56242 6244 56252
rect 6860 56242 6916 56254
rect 7532 56308 7588 56318
rect 7756 56308 7812 59200
rect 7532 56306 7812 56308
rect 7532 56254 7534 56306
rect 7586 56254 7812 56306
rect 7532 56252 7812 56254
rect 8204 56306 8260 59200
rect 8204 56254 8206 56306
rect 8258 56254 8260 56306
rect 7532 56242 7588 56252
rect 8204 56242 8260 56254
rect 8876 56308 8932 56318
rect 9100 56308 9156 59200
rect 8876 56306 9156 56308
rect 8876 56254 8878 56306
rect 8930 56254 9156 56306
rect 8876 56252 9156 56254
rect 8876 56242 8932 56252
rect 5740 55188 5796 55198
rect 5516 55186 5796 55188
rect 5516 55134 5742 55186
rect 5794 55134 5796 55186
rect 5516 55132 5796 55134
rect 9548 55188 9604 59200
rect 10108 56308 10164 56318
rect 10444 56308 10500 59200
rect 10108 56306 10500 56308
rect 10108 56254 10110 56306
rect 10162 56254 10500 56306
rect 10108 56252 10500 56254
rect 10780 56308 10836 56318
rect 10892 56308 10948 59200
rect 10780 56306 10948 56308
rect 10780 56254 10782 56306
rect 10834 56254 10948 56306
rect 10780 56252 10948 56254
rect 10108 56242 10164 56252
rect 10780 56242 10836 56252
rect 11452 56196 11508 56206
rect 11452 56102 11508 56140
rect 11788 56196 11844 59200
rect 12124 56308 12180 56318
rect 12236 56308 12292 59200
rect 12124 56306 12292 56308
rect 12124 56254 12126 56306
rect 12178 56254 12292 56306
rect 12124 56252 12292 56254
rect 12124 56242 12180 56252
rect 11788 56130 11844 56140
rect 12796 55972 12852 55982
rect 13132 55972 13188 59200
rect 12796 55970 13188 55972
rect 12796 55918 12798 55970
rect 12850 55918 13188 55970
rect 12796 55916 13188 55918
rect 12796 55906 12852 55916
rect 9772 55188 9828 55198
rect 9548 55186 9828 55188
rect 9548 55134 9774 55186
rect 9826 55134 9828 55186
rect 9548 55132 9828 55134
rect 13580 55188 13636 59200
rect 14476 57652 14532 59200
rect 14028 57596 14532 57652
rect 14028 55970 14084 57596
rect 14700 56308 14756 56318
rect 14924 56308 14980 59200
rect 15820 57652 15876 59200
rect 14700 56306 14980 56308
rect 14700 56254 14702 56306
rect 14754 56254 14980 56306
rect 14700 56252 14980 56254
rect 15372 57596 15876 57652
rect 14700 56242 14756 56252
rect 14028 55918 14030 55970
rect 14082 55918 14084 55970
rect 14028 55906 14084 55918
rect 15372 55970 15428 57596
rect 16044 56308 16100 56318
rect 16268 56308 16324 59200
rect 16044 56306 16324 56308
rect 16044 56254 16046 56306
rect 16098 56254 16324 56306
rect 16044 56252 16324 56254
rect 16044 56242 16100 56252
rect 15372 55918 15374 55970
rect 15426 55918 15428 55970
rect 15372 55906 15428 55918
rect 16716 55972 16772 55982
rect 16716 55878 16772 55916
rect 17164 55972 17220 59200
rect 17612 56308 17668 59200
rect 17836 56308 17892 56318
rect 17612 56306 17892 56308
rect 17612 56254 17838 56306
rect 17890 56254 17892 56306
rect 17612 56252 17892 56254
rect 17836 56242 17892 56252
rect 17164 55906 17220 55916
rect 18508 55970 18564 59200
rect 18956 56308 19012 59200
rect 19852 57428 19908 59200
rect 19628 57372 19908 57428
rect 19180 56308 19236 56318
rect 18956 56306 19236 56308
rect 18956 56254 19182 56306
rect 19234 56254 19236 56306
rect 18956 56252 19236 56254
rect 19180 56242 19236 56252
rect 18508 55918 18510 55970
rect 18562 55918 18564 55970
rect 18508 55906 18564 55918
rect 19628 55860 19684 57372
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 19964 56308 20020 56318
rect 20300 56308 20356 59200
rect 19964 56306 20356 56308
rect 19964 56254 19966 56306
rect 20018 56254 20356 56306
rect 19964 56252 20356 56254
rect 20636 56642 20692 56654
rect 20636 56590 20638 56642
rect 20690 56590 20692 56642
rect 19964 56242 20020 56252
rect 20636 55970 20692 56590
rect 21196 56642 21252 59200
rect 21196 56590 21198 56642
rect 21250 56590 21252 56642
rect 21196 56578 21252 56590
rect 21644 56308 21700 59200
rect 21756 56308 21812 56318
rect 21644 56306 21812 56308
rect 21644 56254 21758 56306
rect 21810 56254 21812 56306
rect 21644 56252 21812 56254
rect 21756 56242 21812 56252
rect 20636 55918 20638 55970
rect 20690 55918 20692 55970
rect 20636 55906 20692 55918
rect 22540 55970 22596 59200
rect 22988 56308 23044 59200
rect 23100 56308 23156 56318
rect 22988 56306 23156 56308
rect 22988 56254 23102 56306
rect 23154 56254 23156 56306
rect 22988 56252 23156 56254
rect 23100 56242 23156 56252
rect 22540 55918 22542 55970
rect 22594 55918 22596 55970
rect 22540 55906 22596 55918
rect 23884 55970 23940 59200
rect 24332 56308 24388 59200
rect 24444 56308 24500 56318
rect 24332 56306 24500 56308
rect 24332 56254 24446 56306
rect 24498 56254 24500 56306
rect 24332 56252 24500 56254
rect 24444 56242 24500 56252
rect 23884 55918 23886 55970
rect 23938 55918 23940 55970
rect 23884 55906 23940 55918
rect 19628 55804 20132 55860
rect 20076 55522 20132 55804
rect 20076 55470 20078 55522
rect 20130 55470 20132 55522
rect 20076 55458 20132 55470
rect 25228 55524 25284 59200
rect 25676 56306 25732 59200
rect 25676 56254 25678 56306
rect 25730 56254 25732 56306
rect 25676 56242 25732 56254
rect 26460 55972 26516 55982
rect 26572 55972 26628 59200
rect 27020 56306 27076 59200
rect 27020 56254 27022 56306
rect 27074 56254 27076 56306
rect 27020 56242 27076 56254
rect 26460 55970 26628 55972
rect 26460 55918 26462 55970
rect 26514 55918 26628 55970
rect 26460 55916 26628 55918
rect 27804 55972 27860 55982
rect 27916 55972 27972 59200
rect 28364 56306 28420 59200
rect 28364 56254 28366 56306
rect 28418 56254 28420 56306
rect 28364 56242 28420 56254
rect 27804 55970 27972 55972
rect 27804 55918 27806 55970
rect 27858 55918 27972 55970
rect 27804 55916 27972 55918
rect 29260 55970 29316 59200
rect 29708 56308 29764 59200
rect 29932 56308 29988 56318
rect 29708 56306 29988 56308
rect 29708 56254 29934 56306
rect 29986 56254 29988 56306
rect 29708 56252 29988 56254
rect 29932 56242 29988 56252
rect 29260 55918 29262 55970
rect 29314 55918 29316 55970
rect 26460 55906 26516 55916
rect 27804 55906 27860 55916
rect 29260 55906 29316 55918
rect 30604 55970 30660 59200
rect 31052 56308 31108 59200
rect 31276 56308 31332 56318
rect 31052 56306 31332 56308
rect 31052 56254 31278 56306
rect 31330 56254 31332 56306
rect 31052 56252 31332 56254
rect 31276 56242 31332 56252
rect 30604 55918 30606 55970
rect 30658 55918 30660 55970
rect 30604 55906 30660 55918
rect 31948 55972 32004 59200
rect 32396 56642 32452 59200
rect 32396 56590 32398 56642
rect 32450 56590 32452 56642
rect 32396 56578 32452 56590
rect 33180 56642 33236 56654
rect 33180 56590 33182 56642
rect 33234 56590 33236 56642
rect 33180 56306 33236 56590
rect 33180 56254 33182 56306
rect 33234 56254 33236 56306
rect 33180 56242 33236 56254
rect 32172 55972 32228 55982
rect 31948 55970 32228 55972
rect 31948 55918 32174 55970
rect 32226 55918 32228 55970
rect 31948 55916 32228 55918
rect 33292 55972 33348 59200
rect 33740 56642 33796 59200
rect 34636 56754 34692 59200
rect 34636 56702 34638 56754
rect 34690 56702 34692 56754
rect 34636 56690 34692 56702
rect 33740 56590 33742 56642
rect 33794 56590 33796 56642
rect 33740 56578 33796 56590
rect 34524 56642 34580 56654
rect 34524 56590 34526 56642
rect 34578 56590 34580 56642
rect 34524 56306 34580 56590
rect 34524 56254 34526 56306
rect 34578 56254 34580 56306
rect 34524 56242 34580 56254
rect 35084 56196 35140 59200
rect 35980 57090 36036 59200
rect 35980 57038 35982 57090
rect 36034 57038 36036 57090
rect 35980 57026 36036 57038
rect 35196 56754 35252 56766
rect 35196 56702 35198 56754
rect 35250 56702 35252 56754
rect 35196 56306 35252 56702
rect 35196 56254 35198 56306
rect 35250 56254 35252 56306
rect 35196 56242 35252 56254
rect 35084 56130 35140 56140
rect 35868 56196 35924 56206
rect 35868 56102 35924 56140
rect 33852 55972 33908 55982
rect 33292 55970 33908 55972
rect 33292 55918 33854 55970
rect 33906 55918 33908 55970
rect 33292 55916 33908 55918
rect 32172 55906 32228 55916
rect 33852 55906 33908 55916
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 25452 55524 25508 55534
rect 25228 55522 25508 55524
rect 25228 55470 25454 55522
rect 25506 55470 25508 55522
rect 25228 55468 25508 55470
rect 25452 55458 25508 55468
rect 13804 55188 13860 55198
rect 13580 55186 13860 55188
rect 13580 55134 13806 55186
rect 13858 55134 13860 55186
rect 13580 55132 13860 55134
rect 36428 55188 36484 59200
rect 37324 57876 37380 59200
rect 37772 57988 37828 59200
rect 37772 57932 37940 57988
rect 37324 57820 37828 57876
rect 37100 57090 37156 57102
rect 37100 57038 37102 57090
rect 37154 57038 37156 57090
rect 37100 56306 37156 57038
rect 37100 56254 37102 56306
rect 37154 56254 37156 56306
rect 37100 56242 37156 56254
rect 37772 56306 37828 57820
rect 37884 56642 37940 57932
rect 38668 57876 38724 59200
rect 39116 57988 39172 59200
rect 39116 57932 39284 57988
rect 38668 57820 39172 57876
rect 37884 56590 37886 56642
rect 37938 56590 37940 56642
rect 37884 56578 37940 56590
rect 38444 56642 38500 56654
rect 38444 56590 38446 56642
rect 38498 56590 38500 56642
rect 37772 56254 37774 56306
rect 37826 56254 37828 56306
rect 37772 56242 37828 56254
rect 38444 56306 38500 56590
rect 38444 56254 38446 56306
rect 38498 56254 38500 56306
rect 38444 56242 38500 56254
rect 39116 56306 39172 57820
rect 39228 56642 39284 57932
rect 39228 56590 39230 56642
rect 39282 56590 39284 56642
rect 39228 56578 39284 56590
rect 39788 56642 39844 56654
rect 39788 56590 39790 56642
rect 39842 56590 39844 56642
rect 39116 56254 39118 56306
rect 39170 56254 39172 56306
rect 39116 56242 39172 56254
rect 39788 56306 39844 56590
rect 39788 56254 39790 56306
rect 39842 56254 39844 56306
rect 39788 56242 39844 56254
rect 40012 56308 40068 59200
rect 40460 56642 40516 59200
rect 40460 56590 40462 56642
rect 40514 56590 40516 56642
rect 40460 56578 40516 56590
rect 40012 56242 40068 56252
rect 41020 56308 41076 56318
rect 41020 56214 41076 56252
rect 41356 56308 41412 59200
rect 41356 56242 41412 56252
rect 41692 56642 41748 56654
rect 41692 56590 41694 56642
rect 41746 56590 41748 56642
rect 41692 56306 41748 56590
rect 41804 56420 41860 59200
rect 41804 56354 41860 56364
rect 41692 56254 41694 56306
rect 41746 56254 41748 56306
rect 41692 56242 41748 56254
rect 42364 56308 42420 56318
rect 42364 56214 42420 56252
rect 42700 56308 42756 59200
rect 42700 56242 42756 56252
rect 43036 56420 43092 56430
rect 43036 56306 43092 56364
rect 43036 56254 43038 56306
rect 43090 56254 43092 56306
rect 43036 56242 43092 56254
rect 36652 55188 36708 55198
rect 36428 55186 36708 55188
rect 36428 55134 36654 55186
rect 36706 55134 36708 55186
rect 36428 55132 36708 55134
rect 43148 55188 43204 59200
rect 44044 56754 44100 59200
rect 44492 56866 44548 59200
rect 44492 56814 44494 56866
rect 44546 56814 44548 56866
rect 44492 56802 44548 56814
rect 44044 56702 44046 56754
rect 44098 56702 44100 56754
rect 44044 56690 44100 56702
rect 44940 56754 44996 56766
rect 44940 56702 44942 56754
rect 44994 56702 44996 56754
rect 43708 56308 43764 56318
rect 43708 56214 43764 56252
rect 44940 56306 44996 56702
rect 45388 56642 45444 59200
rect 45388 56590 45390 56642
rect 45442 56590 45444 56642
rect 45388 56578 45444 56590
rect 45612 56866 45668 56878
rect 45612 56814 45614 56866
rect 45666 56814 45668 56866
rect 44940 56254 44942 56306
rect 44994 56254 44996 56306
rect 44940 56242 44996 56254
rect 45612 56306 45668 56814
rect 45836 56754 45892 59200
rect 45836 56702 45838 56754
rect 45890 56702 45892 56754
rect 45836 56690 45892 56702
rect 45612 56254 45614 56306
rect 45666 56254 45668 56306
rect 45612 56242 45668 56254
rect 46284 56642 46340 56654
rect 46284 56590 46286 56642
rect 46338 56590 46340 56642
rect 46284 56306 46340 56590
rect 46284 56254 46286 56306
rect 46338 56254 46340 56306
rect 46284 56242 46340 56254
rect 46732 56196 46788 59200
rect 46956 56754 47012 56766
rect 46956 56702 46958 56754
rect 47010 56702 47012 56754
rect 46956 56306 47012 56702
rect 46956 56254 46958 56306
rect 47010 56254 47012 56306
rect 46956 56242 47012 56254
rect 46732 56130 46788 56140
rect 43372 55188 43428 55198
rect 43148 55186 43428 55188
rect 43148 55134 43374 55186
rect 43426 55134 43428 55186
rect 43148 55132 43428 55134
rect 47180 55188 47236 59200
rect 48076 56308 48132 59200
rect 48524 56756 48580 59200
rect 48748 56756 48804 56766
rect 48524 56754 48804 56756
rect 48524 56702 48750 56754
rect 48802 56702 48804 56754
rect 48524 56700 48804 56702
rect 48748 56690 48804 56700
rect 49420 56642 49476 59200
rect 49420 56590 49422 56642
rect 49474 56590 49476 56642
rect 49420 56578 49476 56590
rect 49532 56754 49588 56766
rect 49532 56702 49534 56754
rect 49586 56702 49588 56754
rect 48076 56242 48132 56252
rect 48860 56308 48916 56318
rect 48860 56214 48916 56252
rect 49532 56306 49588 56702
rect 49868 56754 49924 59200
rect 49868 56702 49870 56754
rect 49922 56702 49924 56754
rect 49868 56690 49924 56702
rect 49532 56254 49534 56306
rect 49586 56254 49588 56306
rect 49532 56242 49588 56254
rect 50204 56642 50260 56654
rect 50204 56590 50206 56642
rect 50258 56590 50260 56642
rect 50204 56306 50260 56590
rect 50764 56642 50820 59200
rect 50764 56590 50766 56642
rect 50818 56590 50820 56642
rect 50764 56578 50820 56590
rect 50876 56754 50932 56766
rect 50876 56702 50878 56754
rect 50930 56702 50932 56754
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 50204 56254 50206 56306
rect 50258 56254 50260 56306
rect 50204 56242 50260 56254
rect 50876 56306 50932 56702
rect 50876 56254 50878 56306
rect 50930 56254 50932 56306
rect 50876 56242 50932 56254
rect 47628 56196 47684 56206
rect 47628 56102 47684 56140
rect 47404 55188 47460 55198
rect 47180 55186 47460 55188
rect 47180 55134 47406 55186
rect 47458 55134 47460 55186
rect 47180 55132 47460 55134
rect 51212 55188 51268 59200
rect 51548 56642 51604 56654
rect 51548 56590 51550 56642
rect 51602 56590 51604 56642
rect 51548 56306 51604 56590
rect 52108 56642 52164 59200
rect 52556 56754 52612 59200
rect 52556 56702 52558 56754
rect 52610 56702 52612 56754
rect 52556 56690 52612 56702
rect 53340 56754 53396 56766
rect 53340 56702 53342 56754
rect 53394 56702 53396 56754
rect 52108 56590 52110 56642
rect 52162 56590 52164 56642
rect 52108 56578 52164 56590
rect 52780 56642 52836 56654
rect 52780 56590 52782 56642
rect 52834 56590 52836 56642
rect 51548 56254 51550 56306
rect 51602 56254 51604 56306
rect 51548 56242 51604 56254
rect 52780 56306 52836 56590
rect 52780 56254 52782 56306
rect 52834 56254 52836 56306
rect 52780 56242 52836 56254
rect 53340 56308 53396 56702
rect 53452 56644 53508 59200
rect 53900 56978 53956 59200
rect 53900 56926 53902 56978
rect 53954 56926 53956 56978
rect 53900 56914 53956 56926
rect 54684 56978 54740 56990
rect 54684 56926 54686 56978
rect 54738 56926 54740 56978
rect 53452 56578 53508 56588
rect 54124 56644 54180 56654
rect 53452 56308 53508 56318
rect 53340 56306 53508 56308
rect 53340 56254 53454 56306
rect 53506 56254 53508 56306
rect 53340 56252 53508 56254
rect 53452 56242 53508 56252
rect 54124 56306 54180 56588
rect 54124 56254 54126 56306
rect 54178 56254 54180 56306
rect 54124 56242 54180 56254
rect 54684 56196 54740 56926
rect 54796 56420 54852 59200
rect 54796 56354 54852 56364
rect 54796 56196 54852 56206
rect 54684 56194 54852 56196
rect 54684 56142 54798 56194
rect 54850 56142 54852 56194
rect 54684 56140 54852 56142
rect 54796 56130 54852 56140
rect 51436 55188 51492 55198
rect 51212 55186 51492 55188
rect 51212 55134 51438 55186
rect 51490 55134 51492 55186
rect 51212 55132 51492 55134
rect 55244 55188 55300 59200
rect 55468 56420 55524 56430
rect 55468 56306 55524 56364
rect 55468 56254 55470 56306
rect 55522 56254 55524 56306
rect 55468 56242 55524 56254
rect 55468 55188 55524 55198
rect 55244 55186 55524 55188
rect 55244 55134 55470 55186
rect 55522 55134 55524 55186
rect 55244 55132 55524 55134
rect 5740 55122 5796 55132
rect 9772 55122 9828 55132
rect 13804 55122 13860 55132
rect 36652 55122 36708 55132
rect 43372 55122 43428 55132
rect 47404 55122 47460 55132
rect 51436 55122 51492 55132
rect 55468 55122 55524 55132
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 14896 0 15008 800
rect 44800 0 44912 800
<< via2 >>
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 11452 56194 11508 56196
rect 11452 56142 11454 56194
rect 11454 56142 11506 56194
rect 11506 56142 11508 56194
rect 11452 56140 11508 56142
rect 11788 56140 11844 56196
rect 16716 55970 16772 55972
rect 16716 55918 16718 55970
rect 16718 55918 16770 55970
rect 16770 55918 16772 55970
rect 16716 55916 16772 55918
rect 17164 55916 17220 55972
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 35084 56140 35140 56196
rect 35868 56194 35924 56196
rect 35868 56142 35870 56194
rect 35870 56142 35922 56194
rect 35922 56142 35924 56194
rect 35868 56140 35924 56142
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 40012 56252 40068 56308
rect 41020 56306 41076 56308
rect 41020 56254 41022 56306
rect 41022 56254 41074 56306
rect 41074 56254 41076 56306
rect 41020 56252 41076 56254
rect 41356 56252 41412 56308
rect 41804 56364 41860 56420
rect 42364 56306 42420 56308
rect 42364 56254 42366 56306
rect 42366 56254 42418 56306
rect 42418 56254 42420 56306
rect 42364 56252 42420 56254
rect 42700 56252 42756 56308
rect 43036 56364 43092 56420
rect 43708 56306 43764 56308
rect 43708 56254 43710 56306
rect 43710 56254 43762 56306
rect 43762 56254 43764 56306
rect 43708 56252 43764 56254
rect 46732 56140 46788 56196
rect 48076 56252 48132 56308
rect 48860 56306 48916 56308
rect 48860 56254 48862 56306
rect 48862 56254 48914 56306
rect 48914 56254 48916 56306
rect 48860 56252 48916 56254
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 47628 56194 47684 56196
rect 47628 56142 47630 56194
rect 47630 56142 47682 56194
rect 47682 56142 47684 56194
rect 47628 56140 47684 56142
rect 53452 56588 53508 56644
rect 54124 56588 54180 56644
rect 54796 56364 54852 56420
rect 55468 56364 55524 56420
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 53442 56588 53452 56644
rect 53508 56588 54124 56644
rect 54180 56588 54190 56644
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 41794 56364 41804 56420
rect 41860 56364 43036 56420
rect 43092 56364 43102 56420
rect 54786 56364 54796 56420
rect 54852 56364 55468 56420
rect 55524 56364 55534 56420
rect 40002 56252 40012 56308
rect 40068 56252 41020 56308
rect 41076 56252 41086 56308
rect 41346 56252 41356 56308
rect 41412 56252 42364 56308
rect 42420 56252 42430 56308
rect 42690 56252 42700 56308
rect 42756 56252 43708 56308
rect 43764 56252 43774 56308
rect 48066 56252 48076 56308
rect 48132 56252 48860 56308
rect 48916 56252 48926 56308
rect 11442 56140 11452 56196
rect 11508 56140 11788 56196
rect 11844 56140 11854 56196
rect 35074 56140 35084 56196
rect 35140 56140 35868 56196
rect 35924 56140 35934 56196
rect 46722 56140 46732 56196
rect 46788 56140 47628 56196
rect 47684 56140 47694 56196
rect 16706 55916 16716 55972
rect 16772 55916 17164 55972
rect 17220 55916 17230 55972
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 $PDK_ROOT/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 $PDK_ROOT/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37
timestamp 1669390400
transform 1 0 5488 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1669390400
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72
timestamp 1669390400
transform 1 0 9408 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_107
timestamp 1669390400
transform 1 0 13328 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1669390400
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1669390400
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1669390400
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1669390400
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1669390400
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1669390400
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1669390400
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_422
timestamp 1669390400
transform 1 0 48608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_454
timestamp 1669390400
transform 1 0 52192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_457
timestamp 1669390400
transform 1 0 52528 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1669390400
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_492 $PDK_ROOT/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 56448 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_508
timestamp 1669390400
transform 1 0 58240 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2 $PDK_ROOT/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66 $PDK_ROOT/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1669390400
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1669390400
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1669390400
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_279
timestamp 1669390400
transform 1 0 32592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_350
timestamp 1669390400
transform 1 0 40544 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1669390400
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_421
timestamp 1669390400
transform 1 0 48496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1669390400
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_428
timestamp 1669390400
transform 1 0 49280 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_492
timestamp 1669390400
transform 1 0 56448 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1669390400
transform 1 0 56896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_499 $PDK_ROOT/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 57232 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_507 $PDK_ROOT/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 58128 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1669390400
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1669390400
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1669390400
transform 1 0 28560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_314
timestamp 1669390400
transform 1 0 36512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_385
timestamp 1669390400
transform 1 0 44464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1669390400
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_456
timestamp 1669390400
transform 1 0 52416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1669390400
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_463
timestamp 1669390400
transform 1 0 53200 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_495
timestamp 1669390400
transform 1 0 56784 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_503
timestamp 1669390400
transform 1 0 57680 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_507
timestamp 1669390400
transform 1 0 58128 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1669390400
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1669390400
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1669390400
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1669390400
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1669390400
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1669390400
transform 1 0 40544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1669390400
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_421
timestamp 1669390400
transform 1 0 48496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1669390400
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_428
timestamp 1669390400
transform 1 0 49280 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1669390400
transform 1 0 56448 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1669390400
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_499
timestamp 1669390400
transform 1 0 57232 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_507
timestamp 1669390400
transform 1 0 58128 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1669390400
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1669390400
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1669390400
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1669390400
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1669390400
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1669390400
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1669390400
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1669390400
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_456
timestamp 1669390400
transform 1 0 52416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1669390400
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_463
timestamp 1669390400
transform 1 0 53200 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_495
timestamp 1669390400
transform 1 0 56784 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_503
timestamp 1669390400
transform 1 0 57680 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_507
timestamp 1669390400
transform 1 0 58128 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1669390400
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1669390400
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1669390400
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1669390400
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1669390400
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1669390400
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1669390400
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1669390400
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_421
timestamp 1669390400
transform 1 0 48496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1669390400
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1669390400
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1669390400
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1669390400
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_499
timestamp 1669390400
transform 1 0 57232 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_507
timestamp 1669390400
transform 1 0 58128 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1669390400
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1669390400
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1669390400
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1669390400
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1669390400
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1669390400
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1669390400
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1669390400
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1669390400
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_463
timestamp 1669390400
transform 1 0 53200 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_495
timestamp 1669390400
transform 1 0 56784 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_503
timestamp 1669390400
transform 1 0 57680 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_507
timestamp 1669390400
transform 1 0 58128 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1669390400
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1669390400
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1669390400
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1669390400
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1669390400
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1669390400
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1669390400
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1669390400
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1669390400
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1669390400
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1669390400
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_499
timestamp 1669390400
transform 1 0 57232 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_507
timestamp 1669390400
transform 1 0 58128 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1669390400
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1669390400
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1669390400
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1669390400
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1669390400
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1669390400
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1669390400
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1669390400
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1669390400
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_463
timestamp 1669390400
transform 1 0 53200 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_495
timestamp 1669390400
transform 1 0 56784 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_503
timestamp 1669390400
transform 1 0 57680 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_507
timestamp 1669390400
transform 1 0 58128 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1669390400
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1669390400
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1669390400
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1669390400
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1669390400
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1669390400
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_421
timestamp 1669390400
transform 1 0 48496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1669390400
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1669390400
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1669390400
transform 1 0 56448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1669390400
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_499
timestamp 1669390400
transform 1 0 57232 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_507
timestamp 1669390400
transform 1 0 58128 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1669390400
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1669390400
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1669390400
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1669390400
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1669390400
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1669390400
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1669390400
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1669390400
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_456
timestamp 1669390400
transform 1 0 52416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1669390400
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_463
timestamp 1669390400
transform 1 0 53200 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_495
timestamp 1669390400
transform 1 0 56784 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_503
timestamp 1669390400
transform 1 0 57680 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_507
timestamp 1669390400
transform 1 0 58128 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1669390400
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1669390400
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1669390400
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1669390400
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1669390400
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1669390400
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1669390400
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1669390400
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1669390400
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1669390400
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1669390400
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_499
timestamp 1669390400
transform 1 0 57232 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_507
timestamp 1669390400
transform 1 0 58128 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1669390400
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1669390400
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1669390400
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1669390400
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1669390400
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1669390400
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1669390400
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1669390400
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1669390400
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1669390400
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1669390400
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_463
timestamp 1669390400
transform 1 0 53200 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_495
timestamp 1669390400
transform 1 0 56784 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_503
timestamp 1669390400
transform 1 0 57680 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_507
timestamp 1669390400
transform 1 0 58128 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1669390400
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1669390400
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1669390400
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1669390400
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1669390400
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1669390400
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1669390400
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1669390400
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1669390400
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1669390400
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1669390400
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1669390400
transform 1 0 56448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1669390400
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_499
timestamp 1669390400
transform 1 0 57232 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_507
timestamp 1669390400
transform 1 0 58128 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1669390400
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1669390400
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1669390400
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1669390400
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1669390400
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1669390400
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1669390400
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1669390400
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1669390400
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1669390400
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_463
timestamp 1669390400
transform 1 0 53200 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_495
timestamp 1669390400
transform 1 0 56784 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_503
timestamp 1669390400
transform 1 0 57680 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_507
timestamp 1669390400
transform 1 0 58128 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1669390400
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1669390400
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1669390400
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1669390400
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1669390400
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1669390400
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1669390400
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1669390400
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_428
timestamp 1669390400
transform 1 0 49280 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1669390400
transform 1 0 56448 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1669390400
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_499
timestamp 1669390400
transform 1 0 57232 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_507
timestamp 1669390400
transform 1 0 58128 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1669390400
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1669390400
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1669390400
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1669390400
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1669390400
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1669390400
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_456
timestamp 1669390400
transform 1 0 52416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1669390400
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_463
timestamp 1669390400
transform 1 0 53200 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_495
timestamp 1669390400
transform 1 0 56784 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_503
timestamp 1669390400
transform 1 0 57680 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_507
timestamp 1669390400
transform 1 0 58128 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1669390400
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1669390400
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1669390400
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1669390400
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1669390400
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1669390400
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1669390400
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1669390400
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1669390400
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_428
timestamp 1669390400
transform 1 0 49280 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_492
timestamp 1669390400
transform 1 0 56448 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1669390400
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_499
timestamp 1669390400
transform 1 0 57232 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_507
timestamp 1669390400
transform 1 0 58128 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1669390400
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1669390400
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1669390400
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1669390400
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1669390400
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1669390400
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1669390400
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_456
timestamp 1669390400
transform 1 0 52416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1669390400
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_463
timestamp 1669390400
transform 1 0 53200 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_495
timestamp 1669390400
transform 1 0 56784 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_503
timestamp 1669390400
transform 1 0 57680 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_507
timestamp 1669390400
transform 1 0 58128 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1669390400
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1669390400
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1669390400
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1669390400
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1669390400
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1669390400
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_421
timestamp 1669390400
transform 1 0 48496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1669390400
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_428
timestamp 1669390400
transform 1 0 49280 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1669390400
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1669390400
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_499
timestamp 1669390400
transform 1 0 57232 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_507
timestamp 1669390400
transform 1 0 58128 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1669390400
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1669390400
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1669390400
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1669390400
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1669390400
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1669390400
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1669390400
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1669390400
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_456
timestamp 1669390400
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1669390400
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_463
timestamp 1669390400
transform 1 0 53200 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_495
timestamp 1669390400
transform 1 0 56784 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_503
timestamp 1669390400
transform 1 0 57680 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_507
timestamp 1669390400
transform 1 0 58128 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1669390400
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1669390400
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1669390400
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1669390400
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1669390400
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1669390400
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_421
timestamp 1669390400
transform 1 0 48496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1669390400
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_428
timestamp 1669390400
transform 1 0 49280 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_492
timestamp 1669390400
transform 1 0 56448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1669390400
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_499
timestamp 1669390400
transform 1 0 57232 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_507
timestamp 1669390400
transform 1 0 58128 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1669390400
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1669390400
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1669390400
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1669390400
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1669390400
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1669390400
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1669390400
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1669390400
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1669390400
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1669390400
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1669390400
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_463
timestamp 1669390400
transform 1 0 53200 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_495
timestamp 1669390400
transform 1 0 56784 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_503
timestamp 1669390400
transform 1 0 57680 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_507
timestamp 1669390400
transform 1 0 58128 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_66
timestamp 1669390400
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1669390400
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1669390400
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1669390400
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1669390400
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1669390400
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_421
timestamp 1669390400
transform 1 0 48496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1669390400
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1669390400
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1669390400
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1669390400
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_499
timestamp 1669390400
transform 1 0 57232 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_507
timestamp 1669390400
transform 1 0 58128 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1669390400
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1669390400
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1669390400
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1669390400
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1669390400
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1669390400
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1669390400
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_456
timestamp 1669390400
transform 1 0 52416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1669390400
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_463
timestamp 1669390400
transform 1 0 53200 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_495
timestamp 1669390400
transform 1 0 56784 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_503
timestamp 1669390400
transform 1 0 57680 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_507
timestamp 1669390400
transform 1 0 58128 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_66
timestamp 1669390400
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1669390400
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1669390400
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1669390400
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1669390400
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1669390400
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_421
timestamp 1669390400
transform 1 0 48496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1669390400
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_428
timestamp 1669390400
transform 1 0 49280 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_492
timestamp 1669390400
transform 1 0 56448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1669390400
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_499
timestamp 1669390400
transform 1 0 57232 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_507
timestamp 1669390400
transform 1 0 58128 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1669390400
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1669390400
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1669390400
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1669390400
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1669390400
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1669390400
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_456
timestamp 1669390400
transform 1 0 52416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1669390400
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_463
timestamp 1669390400
transform 1 0 53200 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_495
timestamp 1669390400
transform 1 0 56784 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_503
timestamp 1669390400
transform 1 0 57680 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_507
timestamp 1669390400
transform 1 0 58128 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1669390400
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1669390400
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1669390400
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1669390400
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1669390400
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1669390400
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_421
timestamp 1669390400
transform 1 0 48496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1669390400
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1669390400
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_492
timestamp 1669390400
transform 1 0 56448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1669390400
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_499
timestamp 1669390400
transform 1 0 57232 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_507
timestamp 1669390400
transform 1 0 58128 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1669390400
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1669390400
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1669390400
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1669390400
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1669390400
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1669390400
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1669390400
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1669390400
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_456
timestamp 1669390400
transform 1 0 52416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1669390400
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_463
timestamp 1669390400
transform 1 0 53200 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_495
timestamp 1669390400
transform 1 0 56784 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_503
timestamp 1669390400
transform 1 0 57680 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_507
timestamp 1669390400
transform 1 0 58128 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1669390400
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1669390400
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1669390400
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1669390400
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1669390400
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_421
timestamp 1669390400
transform 1 0 48496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1669390400
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1669390400
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_492
timestamp 1669390400
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1669390400
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_499
timestamp 1669390400
transform 1 0 57232 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_507
timestamp 1669390400
transform 1 0 58128 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1669390400
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1669390400
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1669390400
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1669390400
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1669390400
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1669390400
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1669390400
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_456
timestamp 1669390400
transform 1 0 52416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1669390400
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_463
timestamp 1669390400
transform 1 0 53200 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_495
timestamp 1669390400
transform 1 0 56784 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_503
timestamp 1669390400
transform 1 0 57680 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_507
timestamp 1669390400
transform 1 0 58128 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1669390400
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1669390400
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1669390400
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1669390400
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1669390400
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1669390400
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1669390400
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_421
timestamp 1669390400
transform 1 0 48496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1669390400
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1669390400
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_492
timestamp 1669390400
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1669390400
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_499
timestamp 1669390400
transform 1 0 57232 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_507
timestamp 1669390400
transform 1 0 58128 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1669390400
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1669390400
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1669390400
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1669390400
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1669390400
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1669390400
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1669390400
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1669390400
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_456
timestamp 1669390400
transform 1 0 52416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1669390400
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_463
timestamp 1669390400
transform 1 0 53200 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_495
timestamp 1669390400
transform 1 0 56784 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_503
timestamp 1669390400
transform 1 0 57680 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_507
timestamp 1669390400
transform 1 0 58128 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1669390400
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1669390400
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1669390400
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1669390400
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1669390400
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1669390400
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_421
timestamp 1669390400
transform 1 0 48496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1669390400
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1669390400
transform 1 0 49280 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_492
timestamp 1669390400
transform 1 0 56448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1669390400
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_499
timestamp 1669390400
transform 1 0 57232 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_507
timestamp 1669390400
transform 1 0 58128 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1669390400
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1669390400
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1669390400
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1669390400
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1669390400
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1669390400
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1669390400
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1669390400
transform 1 0 52416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1669390400
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_463
timestamp 1669390400
transform 1 0 53200 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_495
timestamp 1669390400
transform 1 0 56784 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_503
timestamp 1669390400
transform 1 0 57680 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_507
timestamp 1669390400
transform 1 0 58128 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1669390400
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1669390400
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1669390400
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1669390400
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1669390400
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1669390400
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1669390400
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_421
timestamp 1669390400
transform 1 0 48496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1669390400
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1669390400
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1669390400
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1669390400
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_499
timestamp 1669390400
transform 1 0 57232 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_507
timestamp 1669390400
transform 1 0 58128 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1669390400
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1669390400
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1669390400
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1669390400
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1669390400
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1669390400
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1669390400
transform 1 0 52416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1669390400
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_463
timestamp 1669390400
transform 1 0 53200 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_495
timestamp 1669390400
transform 1 0 56784 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_503
timestamp 1669390400
transform 1 0 57680 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_507
timestamp 1669390400
transform 1 0 58128 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1669390400
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1669390400
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1669390400
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1669390400
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1669390400
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1669390400
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1669390400
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_421
timestamp 1669390400
transform 1 0 48496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1669390400
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_428
timestamp 1669390400
transform 1 0 49280 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_492
timestamp 1669390400
transform 1 0 56448 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1669390400
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_499
timestamp 1669390400
transform 1 0 57232 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_507
timestamp 1669390400
transform 1 0 58128 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1669390400
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1669390400
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1669390400
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1669390400
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1669390400
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1669390400
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_456
timestamp 1669390400
transform 1 0 52416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1669390400
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_463
timestamp 1669390400
transform 1 0 53200 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_495
timestamp 1669390400
transform 1 0 56784 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_503
timestamp 1669390400
transform 1 0 57680 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_507
timestamp 1669390400
transform 1 0 58128 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1669390400
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1669390400
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1669390400
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1669390400
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1669390400
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1669390400
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1669390400
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_421
timestamp 1669390400
transform 1 0 48496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1669390400
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1669390400
transform 1 0 49280 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1669390400
transform 1 0 56448 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1669390400
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_499
timestamp 1669390400
transform 1 0 57232 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_507
timestamp 1669390400
transform 1 0 58128 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1669390400
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1669390400
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1669390400
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1669390400
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1669390400
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1669390400
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1669390400
transform 1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1669390400
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_456
timestamp 1669390400
transform 1 0 52416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1669390400
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_463
timestamp 1669390400
transform 1 0 53200 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_495
timestamp 1669390400
transform 1 0 56784 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_503
timestamp 1669390400
transform 1 0 57680 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_507
timestamp 1669390400
transform 1 0 58128 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1669390400
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1669390400
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1669390400
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1669390400
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1669390400
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1669390400
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1669390400
transform 1 0 40544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_421
timestamp 1669390400
transform 1 0 48496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1669390400
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_428
timestamp 1669390400
transform 1 0 49280 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_492
timestamp 1669390400
transform 1 0 56448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1669390400
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_499
timestamp 1669390400
transform 1 0 57232 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_507
timestamp 1669390400
transform 1 0 58128 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1669390400
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1669390400
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_108
timestamp 1669390400
transform 1 0 13440 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_172
timestamp 1669390400
transform 1 0 20608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1669390400
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1669390400
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1669390400
transform 1 0 28560 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_250
timestamp 1669390400
transform 1 0 29344 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_314
timestamp 1669390400
transform 1 0 36512 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1669390400
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_321
timestamp 1669390400
transform 1 0 37296 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_385
timestamp 1669390400
transform 1 0 44464 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1669390400
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_392
timestamp 1669390400
transform 1 0 45248 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_456
timestamp 1669390400
transform 1 0 52416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_460
timestamp 1669390400
transform 1 0 52864 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_463
timestamp 1669390400
transform 1 0 53200 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_495
timestamp 1669390400
transform 1 0 56784 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_503
timestamp 1669390400
transform 1 0 57680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_507
timestamp 1669390400
transform 1 0 58128 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_66
timestamp 1669390400
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1669390400
transform 1 0 9184 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1669390400
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1669390400
transform 1 0 16688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1669390400
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1669390400
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1669390400
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1669390400
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1669390400
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1669390400
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1669390400
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_286
timestamp 1669390400
transform 1 0 33376 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_350
timestamp 1669390400
transform 1 0 40544 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1669390400
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_357
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_421
timestamp 1669390400
transform 1 0 48496 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_425
timestamp 1669390400
transform 1 0 48944 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_428
timestamp 1669390400
transform 1 0 49280 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_492
timestamp 1669390400
transform 1 0 56448 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_496
timestamp 1669390400
transform 1 0 56896 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_499
timestamp 1669390400
transform 1 0 57232 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_507
timestamp 1669390400
transform 1 0 58128 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1669390400
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1669390400
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1669390400
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1669390400
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1669390400
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1669390400
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1669390400
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1669390400
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1669390400
transform 1 0 28560 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1669390400
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1669390400
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1669390400
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1669390400
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_321
timestamp 1669390400
transform 1 0 37296 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1669390400
transform 1 0 44464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1669390400
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_392
timestamp 1669390400
transform 1 0 45248 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_456
timestamp 1669390400
transform 1 0 52416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_460
timestamp 1669390400
transform 1 0 52864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_463
timestamp 1669390400
transform 1 0 53200 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_495
timestamp 1669390400
transform 1 0 56784 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_503
timestamp 1669390400
transform 1 0 57680 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_507
timestamp 1669390400
transform 1 0 58128 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_66
timestamp 1669390400
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1669390400
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1669390400
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1669390400
transform 1 0 16688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1669390400
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1669390400
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1669390400
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1669390400
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1669390400
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1669390400
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1669390400
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1669390400
transform 1 0 33376 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1669390400
transform 1 0 40544 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1669390400
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_357
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_421
timestamp 1669390400
transform 1 0 48496 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_425
timestamp 1669390400
transform 1 0 48944 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_428
timestamp 1669390400
transform 1 0 49280 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_492
timestamp 1669390400
transform 1 0 56448 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_496
timestamp 1669390400
transform 1 0 56896 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_499
timestamp 1669390400
transform 1 0 57232 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_507
timestamp 1669390400
transform 1 0 58128 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1669390400
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1669390400
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1669390400
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1669390400
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1669390400
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1669390400
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1669390400
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1669390400
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1669390400
transform 1 0 28560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1669390400
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1669390400
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1669390400
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1669390400
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_321
timestamp 1669390400
transform 1 0 37296 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_385
timestamp 1669390400
transform 1 0 44464 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1669390400
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_392
timestamp 1669390400
transform 1 0 45248 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_456
timestamp 1669390400
transform 1 0 52416 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_460
timestamp 1669390400
transform 1 0 52864 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_463
timestamp 1669390400
transform 1 0 53200 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_495
timestamp 1669390400
transform 1 0 56784 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_503
timestamp 1669390400
transform 1 0 57680 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_507
timestamp 1669390400
transform 1 0 58128 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_66
timestamp 1669390400
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1669390400
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_73
timestamp 1669390400
transform 1 0 9520 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_137
timestamp 1669390400
transform 1 0 16688 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1669390400
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_144
timestamp 1669390400
transform 1 0 17472 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_208
timestamp 1669390400
transform 1 0 24640 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1669390400
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_215
timestamp 1669390400
transform 1 0 25424 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_279
timestamp 1669390400
transform 1 0 32592 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1669390400
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_286
timestamp 1669390400
transform 1 0 33376 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_350
timestamp 1669390400
transform 1 0 40544 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1669390400
transform 1 0 40992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_357
timestamp 1669390400
transform 1 0 41328 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_421
timestamp 1669390400
transform 1 0 48496 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_425
timestamp 1669390400
transform 1 0 48944 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_428
timestamp 1669390400
transform 1 0 49280 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_492
timestamp 1669390400
transform 1 0 56448 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_496
timestamp 1669390400
transform 1 0 56896 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_499
timestamp 1669390400
transform 1 0 57232 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_507
timestamp 1669390400
transform 1 0 58128 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_2
timestamp 1669390400
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1669390400
transform 1 0 5152 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_37
timestamp 1669390400
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_101
timestamp 1669390400
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1669390400
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_108
timestamp 1669390400
transform 1 0 13440 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_172
timestamp 1669390400
transform 1 0 20608 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1669390400
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_179
timestamp 1669390400
transform 1 0 21392 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_243
timestamp 1669390400
transform 1 0 28560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1669390400
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1669390400
transform 1 0 29344 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_314
timestamp 1669390400
transform 1 0 36512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1669390400
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_321
timestamp 1669390400
transform 1 0 37296 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_385
timestamp 1669390400
transform 1 0 44464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1669390400
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_392
timestamp 1669390400
transform 1 0 45248 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_456
timestamp 1669390400
transform 1 0 52416 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_460
timestamp 1669390400
transform 1 0 52864 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_463
timestamp 1669390400
transform 1 0 53200 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_495
timestamp 1669390400
transform 1 0 56784 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_503
timestamp 1669390400
transform 1 0 57680 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_507
timestamp 1669390400
transform 1 0 58128 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_2
timestamp 1669390400
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_66
timestamp 1669390400
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1669390400
transform 1 0 9184 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_73
timestamp 1669390400
transform 1 0 9520 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_137
timestamp 1669390400
transform 1 0 16688 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1669390400
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_144
timestamp 1669390400
transform 1 0 17472 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_208
timestamp 1669390400
transform 1 0 24640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1669390400
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1669390400
transform 1 0 25424 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1669390400
transform 1 0 32592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1669390400
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1669390400
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1669390400
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1669390400
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_357
timestamp 1669390400
transform 1 0 41328 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_421
timestamp 1669390400
transform 1 0 48496 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_425
timestamp 1669390400
transform 1 0 48944 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_428
timestamp 1669390400
transform 1 0 49280 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_492
timestamp 1669390400
transform 1 0 56448 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_496
timestamp 1669390400
transform 1 0 56896 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_499
timestamp 1669390400
transform 1 0 57232 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_507
timestamp 1669390400
transform 1 0 58128 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_2
timestamp 1669390400
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1669390400
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_37
timestamp 1669390400
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_101
timestamp 1669390400
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1669390400
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_108
timestamp 1669390400
transform 1 0 13440 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_172
timestamp 1669390400
transform 1 0 20608 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1669390400
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1669390400
transform 1 0 21392 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_243
timestamp 1669390400
transform 1 0 28560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1669390400
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_250
timestamp 1669390400
transform 1 0 29344 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_314
timestamp 1669390400
transform 1 0 36512 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1669390400
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_321
timestamp 1669390400
transform 1 0 37296 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_385
timestamp 1669390400
transform 1 0 44464 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1669390400
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_392
timestamp 1669390400
transform 1 0 45248 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_456
timestamp 1669390400
transform 1 0 52416 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_460
timestamp 1669390400
transform 1 0 52864 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_463
timestamp 1669390400
transform 1 0 53200 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_495
timestamp 1669390400
transform 1 0 56784 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_503
timestamp 1669390400
transform 1 0 57680 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_507
timestamp 1669390400
transform 1 0 58128 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_2
timestamp 1669390400
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_66
timestamp 1669390400
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1669390400
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_73
timestamp 1669390400
transform 1 0 9520 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_137
timestamp 1669390400
transform 1 0 16688 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1669390400
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_144
timestamp 1669390400
transform 1 0 17472 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_208
timestamp 1669390400
transform 1 0 24640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1669390400
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_215
timestamp 1669390400
transform 1 0 25424 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_279
timestamp 1669390400
transform 1 0 32592 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1669390400
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1669390400
transform 1 0 33376 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_350
timestamp 1669390400
transform 1 0 40544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1669390400
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_357
timestamp 1669390400
transform 1 0 41328 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_421
timestamp 1669390400
transform 1 0 48496 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_425
timestamp 1669390400
transform 1 0 48944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_428
timestamp 1669390400
transform 1 0 49280 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_492
timestamp 1669390400
transform 1 0 56448 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_496
timestamp 1669390400
transform 1 0 56896 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_499
timestamp 1669390400
transform 1 0 57232 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_507
timestamp 1669390400
transform 1 0 58128 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_2
timestamp 1669390400
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1669390400
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1669390400
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1669390400
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1669390400
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_108
timestamp 1669390400
transform 1 0 13440 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_172
timestamp 1669390400
transform 1 0 20608 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1669390400
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1669390400
transform 1 0 21392 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_243
timestamp 1669390400
transform 1 0 28560 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1669390400
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_250
timestamp 1669390400
transform 1 0 29344 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_314
timestamp 1669390400
transform 1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1669390400
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_321
timestamp 1669390400
transform 1 0 37296 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_385
timestamp 1669390400
transform 1 0 44464 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1669390400
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_392
timestamp 1669390400
transform 1 0 45248 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_456
timestamp 1669390400
transform 1 0 52416 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_460
timestamp 1669390400
transform 1 0 52864 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_463
timestamp 1669390400
transform 1 0 53200 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_495
timestamp 1669390400
transform 1 0 56784 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_503
timestamp 1669390400
transform 1 0 57680 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_507
timestamp 1669390400
transform 1 0 58128 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_2
timestamp 1669390400
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_66
timestamp 1669390400
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1669390400
transform 1 0 9184 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_73
timestamp 1669390400
transform 1 0 9520 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_137
timestamp 1669390400
transform 1 0 16688 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1669390400
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_144
timestamp 1669390400
transform 1 0 17472 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_208
timestamp 1669390400
transform 1 0 24640 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1669390400
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_215
timestamp 1669390400
transform 1 0 25424 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_279
timestamp 1669390400
transform 1 0 32592 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1669390400
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_286
timestamp 1669390400
transform 1 0 33376 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_350
timestamp 1669390400
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1669390400
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_357
timestamp 1669390400
transform 1 0 41328 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_421
timestamp 1669390400
transform 1 0 48496 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_425
timestamp 1669390400
transform 1 0 48944 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_428
timestamp 1669390400
transform 1 0 49280 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_492
timestamp 1669390400
transform 1 0 56448 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_496
timestamp 1669390400
transform 1 0 56896 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_499
timestamp 1669390400
transform 1 0 57232 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_507
timestamp 1669390400
transform 1 0 58128 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_2
timestamp 1669390400
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1669390400
transform 1 0 5152 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_37
timestamp 1669390400
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_101
timestamp 1669390400
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1669390400
transform 1 0 13104 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_108
timestamp 1669390400
transform 1 0 13440 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_172
timestamp 1669390400
transform 1 0 20608 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_176
timestamp 1669390400
transform 1 0 21056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_179
timestamp 1669390400
transform 1 0 21392 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_243
timestamp 1669390400
transform 1 0 28560 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1669390400
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_250
timestamp 1669390400
transform 1 0 29344 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_314
timestamp 1669390400
transform 1 0 36512 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_318
timestamp 1669390400
transform 1 0 36960 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_321
timestamp 1669390400
transform 1 0 37296 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_385
timestamp 1669390400
transform 1 0 44464 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_389
timestamp 1669390400
transform 1 0 44912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_392
timestamp 1669390400
transform 1 0 45248 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_456
timestamp 1669390400
transform 1 0 52416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_460
timestamp 1669390400
transform 1 0 52864 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_463
timestamp 1669390400
transform 1 0 53200 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_495
timestamp 1669390400
transform 1 0 56784 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_503
timestamp 1669390400
transform 1 0 57680 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_507
timestamp 1669390400
transform 1 0 58128 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_2
timestamp 1669390400
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_66
timestamp 1669390400
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_70
timestamp 1669390400
transform 1 0 9184 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_73
timestamp 1669390400
transform 1 0 9520 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_137
timestamp 1669390400
transform 1 0 16688 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_141
timestamp 1669390400
transform 1 0 17136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_144
timestamp 1669390400
transform 1 0 17472 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_208
timestamp 1669390400
transform 1 0 24640 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1669390400
transform 1 0 25088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_215
timestamp 1669390400
transform 1 0 25424 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_279
timestamp 1669390400
transform 1 0 32592 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1669390400
transform 1 0 33040 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_286
timestamp 1669390400
transform 1 0 33376 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_350
timestamp 1669390400
transform 1 0 40544 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1669390400
transform 1 0 40992 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_357
timestamp 1669390400
transform 1 0 41328 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_421
timestamp 1669390400
transform 1 0 48496 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_425
timestamp 1669390400
transform 1 0 48944 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_428
timestamp 1669390400
transform 1 0 49280 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_492
timestamp 1669390400
transform 1 0 56448 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_496
timestamp 1669390400
transform 1 0 56896 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_499
timestamp 1669390400
transform 1 0 57232 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_507
timestamp 1669390400
transform 1 0 58128 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_2
timestamp 1669390400
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1669390400
transform 1 0 5152 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_37
timestamp 1669390400
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_101
timestamp 1669390400
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1669390400
transform 1 0 13104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_108
timestamp 1669390400
transform 1 0 13440 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_172
timestamp 1669390400
transform 1 0 20608 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_176
timestamp 1669390400
transform 1 0 21056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_179
timestamp 1669390400
transform 1 0 21392 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_243
timestamp 1669390400
transform 1 0 28560 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_247
timestamp 1669390400
transform 1 0 29008 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_250
timestamp 1669390400
transform 1 0 29344 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_314
timestamp 1669390400
transform 1 0 36512 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_318
timestamp 1669390400
transform 1 0 36960 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_321
timestamp 1669390400
transform 1 0 37296 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_385
timestamp 1669390400
transform 1 0 44464 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_389
timestamp 1669390400
transform 1 0 44912 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_392
timestamp 1669390400
transform 1 0 45248 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_456
timestamp 1669390400
transform 1 0 52416 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_460
timestamp 1669390400
transform 1 0 52864 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_463
timestamp 1669390400
transform 1 0 53200 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_495
timestamp 1669390400
transform 1 0 56784 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_503
timestamp 1669390400
transform 1 0 57680 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_507
timestamp 1669390400
transform 1 0 58128 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_2
timestamp 1669390400
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_66
timestamp 1669390400
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_70
timestamp 1669390400
transform 1 0 9184 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_73
timestamp 1669390400
transform 1 0 9520 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_137
timestamp 1669390400
transform 1 0 16688 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_141
timestamp 1669390400
transform 1 0 17136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_144
timestamp 1669390400
transform 1 0 17472 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_208
timestamp 1669390400
transform 1 0 24640 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1669390400
transform 1 0 25088 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_215
timestamp 1669390400
transform 1 0 25424 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_279
timestamp 1669390400
transform 1 0 32592 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_283
timestamp 1669390400
transform 1 0 33040 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_286
timestamp 1669390400
transform 1 0 33376 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_350
timestamp 1669390400
transform 1 0 40544 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_354
timestamp 1669390400
transform 1 0 40992 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_357
timestamp 1669390400
transform 1 0 41328 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_421
timestamp 1669390400
transform 1 0 48496 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_425
timestamp 1669390400
transform 1 0 48944 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_428
timestamp 1669390400
transform 1 0 49280 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_492
timestamp 1669390400
transform 1 0 56448 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_496
timestamp 1669390400
transform 1 0 56896 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_499
timestamp 1669390400
transform 1 0 57232 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_507
timestamp 1669390400
transform 1 0 58128 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_2
timestamp 1669390400
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1669390400
transform 1 0 5152 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_37
timestamp 1669390400
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_101
timestamp 1669390400
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1669390400
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_108
timestamp 1669390400
transform 1 0 13440 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_172
timestamp 1669390400
transform 1 0 20608 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_176
timestamp 1669390400
transform 1 0 21056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_179
timestamp 1669390400
transform 1 0 21392 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_243
timestamp 1669390400
transform 1 0 28560 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_247
timestamp 1669390400
transform 1 0 29008 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_250
timestamp 1669390400
transform 1 0 29344 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_314
timestamp 1669390400
transform 1 0 36512 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_318
timestamp 1669390400
transform 1 0 36960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_321
timestamp 1669390400
transform 1 0 37296 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_385
timestamp 1669390400
transform 1 0 44464 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_389
timestamp 1669390400
transform 1 0 44912 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_392
timestamp 1669390400
transform 1 0 45248 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_456
timestamp 1669390400
transform 1 0 52416 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_460
timestamp 1669390400
transform 1 0 52864 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_463
timestamp 1669390400
transform 1 0 53200 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_495
timestamp 1669390400
transform 1 0 56784 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_503
timestamp 1669390400
transform 1 0 57680 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_507
timestamp 1669390400
transform 1 0 58128 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_2
timestamp 1669390400
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_66
timestamp 1669390400
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_70
timestamp 1669390400
transform 1 0 9184 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_73
timestamp 1669390400
transform 1 0 9520 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_137
timestamp 1669390400
transform 1 0 16688 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_141
timestamp 1669390400
transform 1 0 17136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_144
timestamp 1669390400
transform 1 0 17472 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_208
timestamp 1669390400
transform 1 0 24640 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1669390400
transform 1 0 25088 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_215
timestamp 1669390400
transform 1 0 25424 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_279
timestamp 1669390400
transform 1 0 32592 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_283
timestamp 1669390400
transform 1 0 33040 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_286
timestamp 1669390400
transform 1 0 33376 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_350
timestamp 1669390400
transform 1 0 40544 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_354
timestamp 1669390400
transform 1 0 40992 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_357
timestamp 1669390400
transform 1 0 41328 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_421
timestamp 1669390400
transform 1 0 48496 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_425
timestamp 1669390400
transform 1 0 48944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_428
timestamp 1669390400
transform 1 0 49280 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_492
timestamp 1669390400
transform 1 0 56448 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_496
timestamp 1669390400
transform 1 0 56896 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_499
timestamp 1669390400
transform 1 0 57232 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_507
timestamp 1669390400
transform 1 0 58128 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_2
timestamp 1669390400
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1669390400
transform 1 0 5152 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_37
timestamp 1669390400
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_101
timestamp 1669390400
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1669390400
transform 1 0 13104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_108
timestamp 1669390400
transform 1 0 13440 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_172
timestamp 1669390400
transform 1 0 20608 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_176
timestamp 1669390400
transform 1 0 21056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_179
timestamp 1669390400
transform 1 0 21392 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_243
timestamp 1669390400
transform 1 0 28560 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1669390400
transform 1 0 29008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_250
timestamp 1669390400
transform 1 0 29344 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_314
timestamp 1669390400
transform 1 0 36512 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1669390400
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_321
timestamp 1669390400
transform 1 0 37296 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_385
timestamp 1669390400
transform 1 0 44464 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1669390400
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_392
timestamp 1669390400
transform 1 0 45248 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_456
timestamp 1669390400
transform 1 0 52416 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_460
timestamp 1669390400
transform 1 0 52864 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_463
timestamp 1669390400
transform 1 0 53200 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_495
timestamp 1669390400
transform 1 0 56784 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_503
timestamp 1669390400
transform 1 0 57680 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_507
timestamp 1669390400
transform 1 0 58128 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_2
timestamp 1669390400
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_66
timestamp 1669390400
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_70
timestamp 1669390400
transform 1 0 9184 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_73
timestamp 1669390400
transform 1 0 9520 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_137
timestamp 1669390400
transform 1 0 16688 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1669390400
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_144
timestamp 1669390400
transform 1 0 17472 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_208
timestamp 1669390400
transform 1 0 24640 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1669390400
transform 1 0 25088 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_215
timestamp 1669390400
transform 1 0 25424 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_279
timestamp 1669390400
transform 1 0 32592 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1669390400
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_286
timestamp 1669390400
transform 1 0 33376 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_350
timestamp 1669390400
transform 1 0 40544 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_354
timestamp 1669390400
transform 1 0 40992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_357
timestamp 1669390400
transform 1 0 41328 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_421
timestamp 1669390400
transform 1 0 48496 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_425
timestamp 1669390400
transform 1 0 48944 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_428
timestamp 1669390400
transform 1 0 49280 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_492
timestamp 1669390400
transform 1 0 56448 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_496
timestamp 1669390400
transform 1 0 56896 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_499
timestamp 1669390400
transform 1 0 57232 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_507
timestamp 1669390400
transform 1 0 58128 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_2
timestamp 1669390400
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1669390400
transform 1 0 5152 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1669390400
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_101
timestamp 1669390400
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1669390400
transform 1 0 13104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_108
timestamp 1669390400
transform 1 0 13440 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_172
timestamp 1669390400
transform 1 0 20608 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_176
timestamp 1669390400
transform 1 0 21056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_179
timestamp 1669390400
transform 1 0 21392 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_243
timestamp 1669390400
transform 1 0 28560 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_247
timestamp 1669390400
transform 1 0 29008 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_250
timestamp 1669390400
transform 1 0 29344 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_314
timestamp 1669390400
transform 1 0 36512 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1669390400
transform 1 0 36960 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_321
timestamp 1669390400
transform 1 0 37296 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_385
timestamp 1669390400
transform 1 0 44464 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1669390400
transform 1 0 44912 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_392
timestamp 1669390400
transform 1 0 45248 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_456
timestamp 1669390400
transform 1 0 52416 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_460
timestamp 1669390400
transform 1 0 52864 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_463
timestamp 1669390400
transform 1 0 53200 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_495
timestamp 1669390400
transform 1 0 56784 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_503
timestamp 1669390400
transform 1 0 57680 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_507
timestamp 1669390400
transform 1 0 58128 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_2
timestamp 1669390400
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_66
timestamp 1669390400
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_70
timestamp 1669390400
transform 1 0 9184 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_73
timestamp 1669390400
transform 1 0 9520 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_137
timestamp 1669390400
transform 1 0 16688 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1669390400
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_144
timestamp 1669390400
transform 1 0 17472 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_208
timestamp 1669390400
transform 1 0 24640 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1669390400
transform 1 0 25088 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_215
timestamp 1669390400
transform 1 0 25424 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_279
timestamp 1669390400
transform 1 0 32592 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1669390400
transform 1 0 33040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_286
timestamp 1669390400
transform 1 0 33376 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_350
timestamp 1669390400
transform 1 0 40544 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1669390400
transform 1 0 40992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_357
timestamp 1669390400
transform 1 0 41328 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_421
timestamp 1669390400
transform 1 0 48496 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_425
timestamp 1669390400
transform 1 0 48944 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_428
timestamp 1669390400
transform 1 0 49280 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_492
timestamp 1669390400
transform 1 0 56448 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_496
timestamp 1669390400
transform 1 0 56896 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_499
timestamp 1669390400
transform 1 0 57232 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_507
timestamp 1669390400
transform 1 0 58128 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_2
timestamp 1669390400
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1669390400
transform 1 0 5152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1669390400
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1669390400
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1669390400
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_108
timestamp 1669390400
transform 1 0 13440 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_172
timestamp 1669390400
transform 1 0 20608 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_176
timestamp 1669390400
transform 1 0 21056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_179
timestamp 1669390400
transform 1 0 21392 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_243
timestamp 1669390400
transform 1 0 28560 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1669390400
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_250
timestamp 1669390400
transform 1 0 29344 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_314
timestamp 1669390400
transform 1 0 36512 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1669390400
transform 1 0 36960 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_321
timestamp 1669390400
transform 1 0 37296 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_385
timestamp 1669390400
transform 1 0 44464 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1669390400
transform 1 0 44912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_392
timestamp 1669390400
transform 1 0 45248 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_456
timestamp 1669390400
transform 1 0 52416 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_460
timestamp 1669390400
transform 1 0 52864 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_463
timestamp 1669390400
transform 1 0 53200 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_495
timestamp 1669390400
transform 1 0 56784 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_503
timestamp 1669390400
transform 1 0 57680 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_507
timestamp 1669390400
transform 1 0 58128 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_2
timestamp 1669390400
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_66
timestamp 1669390400
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_70
timestamp 1669390400
transform 1 0 9184 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_73
timestamp 1669390400
transform 1 0 9520 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_137
timestamp 1669390400
transform 1 0 16688 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1669390400
transform 1 0 17136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_144
timestamp 1669390400
transform 1 0 17472 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_208
timestamp 1669390400
transform 1 0 24640 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1669390400
transform 1 0 25088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_215
timestamp 1669390400
transform 1 0 25424 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_279
timestamp 1669390400
transform 1 0 32592 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1669390400
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_286
timestamp 1669390400
transform 1 0 33376 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_350
timestamp 1669390400
transform 1 0 40544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1669390400
transform 1 0 40992 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_357
timestamp 1669390400
transform 1 0 41328 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_421
timestamp 1669390400
transform 1 0 48496 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_425
timestamp 1669390400
transform 1 0 48944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_428
timestamp 1669390400
transform 1 0 49280 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_492
timestamp 1669390400
transform 1 0 56448 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_496
timestamp 1669390400
transform 1 0 56896 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_499
timestamp 1669390400
transform 1 0 57232 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_507
timestamp 1669390400
transform 1 0 58128 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_2
timestamp 1669390400
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_34
timestamp 1669390400
transform 1 0 5152 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_37
timestamp 1669390400
transform 1 0 5488 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_42
timestamp 1669390400
transform 1 0 6048 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_78
timestamp 1669390400
transform 1 0 10080 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_94
timestamp 1669390400
transform 1 0 11872 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_102
timestamp 1669390400
transform 1 0 12768 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_108
timestamp 1669390400
transform 1 0 13440 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_114
timestamp 1669390400
transform 1 0 14112 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_146
timestamp 1669390400
transform 1 0 17696 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_162
timestamp 1669390400
transform 1 0 19488 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_170
timestamp 1669390400
transform 1 0 20384 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_174
timestamp 1669390400
transform 1 0 20832 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_176
timestamp 1669390400
transform 1 0 21056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_179
timestamp 1669390400
transform 1 0 21392 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_211
timestamp 1669390400
transform 1 0 24976 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_213
timestamp 1669390400
transform 1 0 25200 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_218
timestamp 1669390400
transform 1 0 25760 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_234
timestamp 1669390400
transform 1 0 27552 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_242
timestamp 1669390400
transform 1 0 28448 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_246
timestamp 1669390400
transform 1 0 28896 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_250
timestamp 1669390400
transform 1 0 29344 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1669390400
transform 1 0 36960 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_321
timestamp 1669390400
transform 1 0 37296 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_353
timestamp 1669390400
transform 1 0 40880 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_369
timestamp 1669390400
transform 1 0 42672 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_373
timestamp 1669390400
transform 1 0 43120 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_378
timestamp 1669390400
transform 1 0 43680 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_386
timestamp 1669390400
transform 1 0 44576 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_392
timestamp 1669390400
transform 1 0 45248 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_408
timestamp 1669390400
transform 1 0 47040 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_414
timestamp 1669390400
transform 1 0 47712 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_450
timestamp 1669390400
transform 1 0 51744 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_458
timestamp 1669390400
transform 1 0 52640 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_460
timestamp 1669390400
transform 1 0 52864 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_463
timestamp 1669390400
transform 1 0 53200 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_479
timestamp 1669390400
transform 1 0 54992 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_481
timestamp 1669390400
transform 1 0 55216 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_486
timestamp 1669390400
transform 1 0 55776 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_502
timestamp 1669390400
transform 1 0 57568 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_506
timestamp 1669390400
transform 1 0 58016 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_508
timestamp 1669390400
transform 1 0 58240 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_2
timestamp 1669390400
transform 1 0 1568 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_18
timestamp 1669390400
transform 1 0 3360 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_26
timestamp 1669390400
transform 1 0 4256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_34
timestamp 1669390400
transform 1 0 5152 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_37
timestamp 1669390400
transform 1 0 5488 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_45
timestamp 1669390400
transform 1 0 6384 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_51
timestamp 1669390400
transform 1 0 7056 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_57
timestamp 1669390400
transform 1 0 7728 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_63
timestamp 1669390400
transform 1 0 8400 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_69
timestamp 1669390400
transform 1 0 9072 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_72
timestamp 1669390400
transform 1 0 9408 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_80
timestamp 1669390400
transform 1 0 10304 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_86
timestamp 1669390400
transform 1 0 10976 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_92
timestamp 1669390400
transform 1 0 11648 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_98
timestamp 1669390400
transform 1 0 12320 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_104
timestamp 1669390400
transform 1 0 12992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_107
timestamp 1669390400
transform 1 0 13328 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_115
timestamp 1669390400
transform 1 0 14224 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_121
timestamp 1669390400
transform 1 0 14896 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_127
timestamp 1669390400
transform 1 0 15568 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_133
timestamp 1669390400
transform 1 0 16240 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_139
timestamp 1669390400
transform 1 0 16912 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_142
timestamp 1669390400
transform 1 0 17248 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_150
timestamp 1669390400
transform 1 0 18144 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_156
timestamp 1669390400
transform 1 0 18816 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_162
timestamp 1669390400
transform 1 0 19488 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_168
timestamp 1669390400
transform 1 0 20160 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_174
timestamp 1669390400
transform 1 0 20832 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_177
timestamp 1669390400
transform 1 0 21168 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_185
timestamp 1669390400
transform 1 0 22064 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_191
timestamp 1669390400
transform 1 0 22736 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_197
timestamp 1669390400
transform 1 0 23408 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_203
timestamp 1669390400
transform 1 0 24080 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_209
timestamp 1669390400
transform 1 0 24752 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_212
timestamp 1669390400
transform 1 0 25088 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_220
timestamp 1669390400
transform 1 0 25984 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_226
timestamp 1669390400
transform 1 0 26656 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_232
timestamp 1669390400
transform 1 0 27328 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_238
timestamp 1669390400
transform 1 0 28000 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_244
timestamp 1669390400
transform 1 0 28672 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_247
timestamp 1669390400
transform 1 0 29008 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_252
timestamp 1669390400
transform 1 0 29568 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_258
timestamp 1669390400
transform 1 0 30240 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_264
timestamp 1669390400
transform 1 0 30912 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_270
timestamp 1669390400
transform 1 0 31584 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_278
timestamp 1669390400
transform 1 0 32480 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_282
timestamp 1669390400
transform 1 0 32928 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_287
timestamp 1669390400
transform 1 0 33488 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_293
timestamp 1669390400
transform 1 0 34160 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_299
timestamp 1669390400
transform 1 0 34832 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_305
timestamp 1669390400
transform 1 0 35504 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_311
timestamp 1669390400
transform 1 0 36176 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_317
timestamp 1669390400
transform 1 0 36848 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_322
timestamp 1669390400
transform 1 0 37408 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_328
timestamp 1669390400
transform 1 0 38080 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_334
timestamp 1669390400
transform 1 0 38752 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_340
timestamp 1669390400
transform 1 0 39424 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_346
timestamp 1669390400
transform 1 0 40096 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_352
timestamp 1669390400
transform 1 0 40768 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_357
timestamp 1669390400
transform 1 0 41328 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_363
timestamp 1669390400
transform 1 0 42000 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_369
timestamp 1669390400
transform 1 0 42672 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_375
timestamp 1669390400
transform 1 0 43344 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_381
timestamp 1669390400
transform 1 0 44016 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_387
timestamp 1669390400
transform 1 0 44688 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_392
timestamp 1669390400
transform 1 0 45248 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_398
timestamp 1669390400
transform 1 0 45920 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_404
timestamp 1669390400
transform 1 0 46592 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_410
timestamp 1669390400
transform 1 0 47264 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_416
timestamp 1669390400
transform 1 0 47936 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_422
timestamp 1669390400
transform 1 0 48608 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_427
timestamp 1669390400
transform 1 0 49168 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_433
timestamp 1669390400
transform 1 0 49840 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_439
timestamp 1669390400
transform 1 0 50512 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_445
timestamp 1669390400
transform 1 0 51184 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_451
timestamp 1669390400
transform 1 0 51856 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_457
timestamp 1669390400
transform 1 0 52528 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_462
timestamp 1669390400
transform 1 0 53088 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_468
timestamp 1669390400
transform 1 0 53760 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_474
timestamp 1669390400
transform 1 0 54432 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_480
timestamp 1669390400
transform 1 0 55104 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_486
timestamp 1669390400
transform 1 0 55776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_492
timestamp 1669390400
transform 1 0 56448 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_508
timestamp 1669390400
transform 1 0 58240 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 $PDK_ROOT/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1669390400
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1669390400
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1669390400
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1669390400
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1669390400
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1669390400
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1669390400
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1669390400
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1669390400
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1669390400
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1669390400
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1669390400
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1669390400
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1669390400
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1669390400
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1669390400
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1669390400
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1669390400
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1669390400
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1669390400
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1669390400
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1669390400
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1669390400
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1669390400
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1669390400
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1669390400
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1669390400
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1669390400
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1669390400
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1669390400
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1669390400
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1669390400
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1669390400
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1669390400
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1669390400
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1669390400
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1669390400
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1669390400
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1669390400
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1669390400
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136 $PDK_ROOT/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1669390400
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1669390400
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1669390400
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1669390400
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1669390400
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1669390400
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1669390400
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1669390400
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1669390400
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1669390400
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1669390400
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1669390400
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1669390400
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1669390400
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1669390400
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1669390400
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1669390400
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1669390400
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1669390400
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1669390400
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1669390400
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1669390400
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1669390400
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1669390400
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1669390400
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1669390400
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1669390400
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1669390400
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1669390400
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1669390400
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1669390400
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1669390400
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1669390400
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1669390400
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1669390400
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1669390400
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1669390400
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1669390400
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1669390400
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1669390400
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1669390400
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1669390400
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1669390400
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1669390400
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1669390400
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1669390400
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1669390400
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1669390400
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1669390400
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1669390400
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1669390400
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1669390400
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1669390400
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1669390400
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1669390400
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1669390400
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1669390400
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1669390400
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1669390400
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1669390400
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1669390400
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1669390400
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1669390400
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1669390400
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1669390400
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1669390400
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1669390400
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1669390400
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1669390400
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1669390400
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1669390400
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1669390400
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1669390400
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1669390400
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1669390400
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1669390400
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1669390400
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1669390400
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1669390400
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1669390400
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1669390400
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1669390400
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1669390400
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1669390400
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1669390400
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1669390400
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1669390400
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1669390400
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1669390400
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1669390400
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1669390400
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1669390400
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1669390400
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1669390400
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1669390400
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1669390400
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1669390400
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1669390400
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1669390400
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1669390400
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1669390400
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1669390400
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1669390400
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1669390400
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1669390400
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1669390400
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1669390400
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1669390400
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1669390400
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1669390400
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1669390400
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1669390400
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1669390400
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1669390400
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1669390400
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1669390400
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1669390400
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1669390400
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1669390400
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1669390400
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1669390400
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1669390400
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1669390400
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1669390400
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1669390400
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1669390400
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1669390400
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1669390400
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1669390400
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1669390400
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1669390400
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1669390400
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1669390400
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1669390400
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1669390400
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1669390400
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1669390400
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1669390400
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1669390400
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1669390400
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1669390400
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1669390400
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1669390400
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1669390400
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1669390400
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1669390400
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1669390400
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1669390400
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1669390400
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1669390400
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1669390400
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1669390400
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1669390400
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1669390400
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1669390400
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1669390400
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1669390400
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1669390400
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1669390400
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1669390400
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1669390400
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1669390400
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1669390400
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1669390400
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1669390400
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1669390400
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1669390400
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1669390400
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1669390400
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1669390400
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1669390400
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1669390400
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1669390400
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1669390400
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1669390400
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1669390400
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1669390400
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1669390400
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1669390400
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1669390400
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1669390400
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1669390400
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1669390400
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1669390400
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1669390400
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1669390400
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1669390400
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1669390400
transform 1 0 5264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1669390400
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1669390400
transform 1 0 13104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1669390400
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1669390400
transform 1 0 20944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1669390400
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1669390400
transform 1 0 28784 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1669390400
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1669390400
transform 1 0 36624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1669390400
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1669390400
transform 1 0 44464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1669390400
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1669390400
transform 1 0 52304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1669390400
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_1 $PDK_ROOT/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4704 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_2
timestamp 1669390400
transform 1 0 5936 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_3
timestamp 1669390400
transform 1 0 7280 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_4
timestamp 1669390400
transform 1 0 8624 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_5
timestamp 1669390400
transform 1 0 9856 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_6
timestamp 1669390400
transform 1 0 11200 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_7
timestamp 1669390400
transform -1 0 35504 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_8
timestamp 1669390400
transform -1 0 37408 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_9
timestamp 1669390400
transform -1 0 38080 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_10
timestamp 1669390400
transform -1 0 39424 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_11
timestamp 1669390400
transform -1 0 41328 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_12
timestamp 1669390400
transform -1 0 42672 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_13
timestamp 1669390400
transform -1 0 44016 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_14
timestamp 1669390400
transform -1 0 45248 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_15
timestamp 1669390400
transform -1 0 46592 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_16
timestamp 1669390400
transform -1 0 47936 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_17
timestamp 1669390400
transform -1 0 49168 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_18
timestamp 1669390400
transform -1 0 50512 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_19
timestamp 1669390400
transform -1 0 51856 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_20
timestamp 1669390400
transform -1 0 53088 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_21
timestamp 1669390400
transform -1 0 54432 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_22
timestamp 1669390400
transform -1 0 55776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_23
timestamp 1669390400
transform -1 0 6048 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_24
timestamp 1669390400
transform 1 0 6608 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_25
timestamp 1669390400
transform 1 0 7952 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_26
timestamp 1669390400
transform -1 0 10080 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_27
timestamp 1669390400
transform 1 0 10528 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_28
timestamp 1669390400
transform 1 0 11872 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_29
timestamp 1669390400
transform -1 0 14112 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_30
timestamp 1669390400
transform 1 0 14448 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_31
timestamp 1669390400
transform 1 0 15792 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_32
timestamp 1669390400
transform -1 0 18144 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_33
timestamp 1669390400
transform -1 0 19488 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_34
timestamp 1669390400
transform 1 0 19712 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_35
timestamp 1669390400
transform -1 0 22064 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_36
timestamp 1669390400
transform -1 0 23408 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_37
timestamp 1669390400
transform -1 0 24752 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_38
timestamp 1669390400
transform -1 0 25984 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_39
timestamp 1669390400
transform -1 0 27328 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_40
timestamp 1669390400
transform -1 0 28672 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_41
timestamp 1669390400
transform -1 0 30240 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_42
timestamp 1669390400
transform -1 0 31584 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_43
timestamp 1669390400
transform -1 0 33488 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_44
timestamp 1669390400
transform -1 0 34832 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_45
timestamp 1669390400
transform -1 0 36176 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_46
timestamp 1669390400
transform -1 0 36960 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_47
timestamp 1669390400
transform -1 0 38752 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_48
timestamp 1669390400
transform -1 0 40096 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_49
timestamp 1669390400
transform -1 0 42000 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_50
timestamp 1669390400
transform -1 0 43344 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_51
timestamp 1669390400
transform -1 0 43680 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_52
timestamp 1669390400
transform -1 0 45920 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_53
timestamp 1669390400
transform -1 0 47264 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_54
timestamp 1669390400
transform -1 0 47712 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_55
timestamp 1669390400
transform -1 0 49840 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_56
timestamp 1669390400
transform -1 0 51184 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_57
timestamp 1669390400
transform -1 0 51744 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_58
timestamp 1669390400
transform -1 0 53760 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_59
timestamp 1669390400
transform -1 0 55104 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_multiplier_8_60
timestamp 1669390400
transform -1 0 55776 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_61 $PDK_ROOT/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 12544 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_62
timestamp 1669390400
transform 1 0 13776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_63
timestamp 1669390400
transform 1 0 15120 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_64
timestamp 1669390400
transform 1 0 16464 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_65
timestamp 1669390400
transform -1 0 18816 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_66
timestamp 1669390400
transform -1 0 20384 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_67
timestamp 1669390400
transform 1 0 20384 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_68
timestamp 1669390400
transform 1 0 22288 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_69
timestamp 1669390400
transform 1 0 23632 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_70
timestamp 1669390400
transform -1 0 25760 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_71
timestamp 1669390400
transform 1 0 26208 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_72
timestamp 1669390400
transform 1 0 27552 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_73
timestamp 1669390400
transform -1 0 29568 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_74
timestamp 1669390400
transform -1 0 30912 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_75
timestamp 1669390400
transform -1 0 32480 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  wrapped_multiplier_8_76
timestamp 1669390400
transform -1 0 34160 0 -1 56448
box -86 -86 534 870
<< labels >>
flabel metal2 s 4592 59200 4704 60000 0 FreeSans 448 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 18032 59200 18144 60000 0 FreeSans 448 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 19376 59200 19488 60000 0 FreeSans 448 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 20720 59200 20832 60000 0 FreeSans 448 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 22064 59200 22176 60000 0 FreeSans 448 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 23408 59200 23520 60000 0 FreeSans 448 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 24752 59200 24864 60000 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 26096 59200 26208 60000 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 27440 59200 27552 60000 0 FreeSans 448 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 28784 59200 28896 60000 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 30128 59200 30240 60000 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal2 s 5936 59200 6048 60000 0 FreeSans 448 90 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 31472 59200 31584 60000 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 32816 59200 32928 60000 0 FreeSans 448 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 34160 59200 34272 60000 0 FreeSans 448 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 35504 59200 35616 60000 0 FreeSans 448 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal2 s 36848 59200 36960 60000 0 FreeSans 448 90 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 38192 59200 38304 60000 0 FreeSans 448 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal2 s 39536 59200 39648 60000 0 FreeSans 448 90 0 0 io_in[26]
port 18 nsew signal input
flabel metal2 s 40880 59200 40992 60000 0 FreeSans 448 90 0 0 io_in[27]
port 19 nsew signal input
flabel metal2 s 42224 59200 42336 60000 0 FreeSans 448 90 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 43568 59200 43680 60000 0 FreeSans 448 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 7280 59200 7392 60000 0 FreeSans 448 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 44912 59200 45024 60000 0 FreeSans 448 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 46256 59200 46368 60000 0 FreeSans 448 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 47600 59200 47712 60000 0 FreeSans 448 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 48944 59200 49056 60000 0 FreeSans 448 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 50288 59200 50400 60000 0 FreeSans 448 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal2 s 51632 59200 51744 60000 0 FreeSans 448 90 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 52976 59200 53088 60000 0 FreeSans 448 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal2 s 54320 59200 54432 60000 0 FreeSans 448 90 0 0 io_in[37]
port 30 nsew signal input
flabel metal2 s 8624 59200 8736 60000 0 FreeSans 448 90 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 9968 59200 10080 60000 0 FreeSans 448 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 11312 59200 11424 60000 0 FreeSans 448 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 12656 59200 12768 60000 0 FreeSans 448 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 14000 59200 14112 60000 0 FreeSans 448 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 15344 59200 15456 60000 0 FreeSans 448 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 16688 59200 16800 60000 0 FreeSans 448 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 5040 59200 5152 60000 0 FreeSans 448 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal2 s 18480 59200 18592 60000 0 FreeSans 448 90 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal2 s 19824 59200 19936 60000 0 FreeSans 448 90 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal2 s 21168 59200 21280 60000 0 FreeSans 448 90 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal2 s 22512 59200 22624 60000 0 FreeSans 448 90 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 23856 59200 23968 60000 0 FreeSans 448 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 25200 59200 25312 60000 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 26544 59200 26656 60000 0 FreeSans 448 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 27888 59200 28000 60000 0 FreeSans 448 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 29232 59200 29344 60000 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 30576 59200 30688 60000 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 6384 59200 6496 60000 0 FreeSans 448 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 31920 59200 32032 60000 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 33264 59200 33376 60000 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 34608 59200 34720 60000 0 FreeSans 448 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 35952 59200 36064 60000 0 FreeSans 448 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal2 s 37296 59200 37408 60000 0 FreeSans 448 90 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 38640 59200 38752 60000 0 FreeSans 448 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 39984 59200 40096 60000 0 FreeSans 448 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal2 s 41328 59200 41440 60000 0 FreeSans 448 90 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal2 s 42672 59200 42784 60000 0 FreeSans 448 90 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal2 s 44016 59200 44128 60000 0 FreeSans 448 90 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 7728 59200 7840 60000 0 FreeSans 448 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 45360 59200 45472 60000 0 FreeSans 448 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal2 s 46704 59200 46816 60000 0 FreeSans 448 90 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal2 s 48048 59200 48160 60000 0 FreeSans 448 90 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal2 s 49392 59200 49504 60000 0 FreeSans 448 90 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal2 s 50736 59200 50848 60000 0 FreeSans 448 90 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal2 s 52080 59200 52192 60000 0 FreeSans 448 90 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 53424 59200 53536 60000 0 FreeSans 448 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal2 s 54768 59200 54880 60000 0 FreeSans 448 90 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal2 s 9072 59200 9184 60000 0 FreeSans 448 90 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 10416 59200 10528 60000 0 FreeSans 448 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal2 s 11760 59200 11872 60000 0 FreeSans 448 90 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal2 s 13104 59200 13216 60000 0 FreeSans 448 90 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal2 s 14448 59200 14560 60000 0 FreeSans 448 90 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal2 s 15792 59200 15904 60000 0 FreeSans 448 90 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 17136 59200 17248 60000 0 FreeSans 448 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal2 s 5488 59200 5600 60000 0 FreeSans 448 90 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 18928 59200 19040 60000 0 FreeSans 448 90 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal2 s 20272 59200 20384 60000 0 FreeSans 448 90 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal2 s 21616 59200 21728 60000 0 FreeSans 448 90 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal2 s 22960 59200 23072 60000 0 FreeSans 448 90 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 24304 59200 24416 60000 0 FreeSans 448 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 25648 59200 25760 60000 0 FreeSans 448 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 26992 59200 27104 60000 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 28336 59200 28448 60000 0 FreeSans 448 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 29680 59200 29792 60000 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 31024 59200 31136 60000 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 6832 59200 6944 60000 0 FreeSans 448 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 32368 59200 32480 60000 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 33712 59200 33824 60000 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 35056 59200 35168 60000 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 36400 59200 36512 60000 0 FreeSans 448 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal2 s 37744 59200 37856 60000 0 FreeSans 448 90 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 39088 59200 39200 60000 0 FreeSans 448 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 40432 59200 40544 60000 0 FreeSans 448 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 41776 59200 41888 60000 0 FreeSans 448 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 43120 59200 43232 60000 0 FreeSans 448 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 44464 59200 44576 60000 0 FreeSans 448 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal2 s 8176 59200 8288 60000 0 FreeSans 448 90 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal2 s 45808 59200 45920 60000 0 FreeSans 448 90 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal2 s 47152 59200 47264 60000 0 FreeSans 448 90 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 48496 59200 48608 60000 0 FreeSans 448 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 49840 59200 49952 60000 0 FreeSans 448 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal2 s 51184 59200 51296 60000 0 FreeSans 448 90 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal2 s 52528 59200 52640 60000 0 FreeSans 448 90 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 53872 59200 53984 60000 0 FreeSans 448 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 55216 59200 55328 60000 0 FreeSans 448 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 9520 59200 9632 60000 0 FreeSans 448 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 10864 59200 10976 60000 0 FreeSans 448 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 12208 59200 12320 60000 0 FreeSans 448 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 13552 59200 13664 60000 0 FreeSans 448 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal2 s 14896 59200 15008 60000 0 FreeSans 448 90 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal2 s 16240 59200 16352 60000 0 FreeSans 448 90 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal2 s 17584 59200 17696 60000 0 FreeSans 448 90 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 114 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 114 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 115 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 115 nsew ground bidirectional
flabel metal2 s 14896 0 15008 800 0 FreeSans 448 90 0 0 wb_clk_i
port 116 nsew signal input
flabel metal2 s 44800 0 44912 800 0 FreeSans 448 90 0 0 wb_rst_i
port 117 nsew signal input
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal2 5040 56280 5040 56280 0 net1
rlabel metal2 39144 57064 39144 57064 0 net10
rlabel metal3 40544 56280 40544 56280 0 net11
rlabel metal3 41888 56280 41888 56280 0 net12
rlabel metal3 43232 56280 43232 56280 0 net13
rlabel metal2 44968 56504 44968 56504 0 net14
rlabel metal2 46312 56448 46312 56448 0 net15
rlabel metal2 46760 57722 46760 57722 0 net16
rlabel metal3 48496 56280 48496 56280 0 net17
rlabel metal2 50232 56448 50232 56448 0 net18
rlabel metal2 51576 56448 51576 56448 0 net19
rlabel metal2 6328 56280 6328 56280 0 net2
rlabel metal2 52808 56448 52808 56448 0 net20
rlabel metal2 54152 56448 54152 56448 0 net21
rlabel metal2 55496 56336 55496 56336 0 net22
rlabel metal2 5656 55160 5656 55160 0 net23
rlabel metal2 6888 57778 6888 57778 0 net24
rlabel metal2 8232 57778 8232 57778 0 net25
rlabel metal2 9688 55160 9688 55160 0 net26
rlabel metal2 10864 56280 10864 56280 0 net27
rlabel metal2 12208 56280 12208 56280 0 net28
rlabel metal2 13720 55160 13720 55160 0 net29
rlabel metal2 7672 56280 7672 56280 0 net3
rlabel metal2 14840 56280 14840 56280 0 net30
rlabel metal2 16184 56280 16184 56280 0 net31
rlabel metal2 17752 56280 17752 56280 0 net32
rlabel metal2 19096 56280 19096 56280 0 net33
rlabel metal2 20160 56280 20160 56280 0 net34
rlabel metal2 21728 56280 21728 56280 0 net35
rlabel metal2 23072 56280 23072 56280 0 net36
rlabel metal2 24416 56280 24416 56280 0 net37
rlabel metal2 25704 57778 25704 57778 0 net38
rlabel metal2 27048 57778 27048 57778 0 net39
rlabel metal2 9016 56280 9016 56280 0 net4
rlabel metal2 28392 57778 28392 57778 0 net40
rlabel metal2 29848 56280 29848 56280 0 net41
rlabel metal2 31192 56280 31192 56280 0 net42
rlabel metal2 33208 56448 33208 56448 0 net43
rlabel metal2 34552 56448 34552 56448 0 net44
rlabel metal2 35112 57722 35112 57722 0 net45
rlabel metal2 36568 55160 36568 55160 0 net46
rlabel metal2 38472 56448 38472 56448 0 net47
rlabel metal2 39816 56448 39816 56448 0 net48
rlabel metal2 41720 56448 41720 56448 0 net49
rlabel metal2 10304 56280 10304 56280 0 net5
rlabel metal2 43064 56336 43064 56336 0 net50
rlabel metal2 43288 55160 43288 55160 0 net51
rlabel metal2 45640 56560 45640 56560 0 net52
rlabel metal2 46984 56504 46984 56504 0 net53
rlabel metal2 47320 55160 47320 55160 0 net54
rlabel metal2 49560 56504 49560 56504 0 net55
rlabel metal2 50904 56504 50904 56504 0 net56
rlabel metal2 51352 55160 51352 55160 0 net57
rlabel metal2 53424 56280 53424 56280 0 net58
rlabel metal2 54768 56168 54768 56168 0 net59
rlabel metal2 11816 57722 11816 57722 0 net6
rlabel metal2 55384 55160 55384 55160 0 net60
rlabel metal2 12992 55944 12992 55944 0 net61
rlabel metal2 14056 56784 14056 56784 0 net62
rlabel metal2 15400 56784 15400 56784 0 net63
rlabel metal3 16968 55944 16968 55944 0 net64
rlabel metal2 18536 57610 18536 57610 0 net65
rlabel metal2 20104 55664 20104 55664 0 net66
rlabel metal2 20664 56280 20664 56280 0 net67
rlabel metal2 22568 57610 22568 57610 0 net68
rlabel metal2 23912 57610 23912 57610 0 net69
rlabel metal2 35224 56504 35224 56504 0 net7
rlabel metal2 25368 55496 25368 55496 0 net70
rlabel metal2 26544 55944 26544 55944 0 net71
rlabel metal2 27888 55944 27888 55944 0 net72
rlabel metal2 29288 57610 29288 57610 0 net73
rlabel metal2 30632 57610 30632 57610 0 net74
rlabel metal2 32088 55944 32088 55944 0 net75
rlabel metal2 33600 55944 33600 55944 0 net76
rlabel metal2 37128 56672 37128 56672 0 net8
rlabel metal2 37800 57064 37800 57064 0 net9
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
