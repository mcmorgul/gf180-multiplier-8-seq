magic
tech gf180mcuC
magscale 1 5
timestamp 1670279682
<< obsm1 >>
rect 672 1538 29288 28545
<< metal2 >>
rect 2296 29600 2352 30000
rect 2520 29600 2576 30000
rect 2744 29600 2800 30000
rect 2968 29600 3024 30000
rect 3192 29600 3248 30000
rect 3416 29600 3472 30000
rect 3640 29600 3696 30000
rect 3864 29600 3920 30000
rect 4088 29600 4144 30000
rect 4312 29600 4368 30000
rect 4536 29600 4592 30000
rect 4760 29600 4816 30000
rect 4984 29600 5040 30000
rect 5208 29600 5264 30000
rect 5432 29600 5488 30000
rect 5656 29600 5712 30000
rect 5880 29600 5936 30000
rect 6104 29600 6160 30000
rect 6328 29600 6384 30000
rect 6552 29600 6608 30000
rect 6776 29600 6832 30000
rect 7000 29600 7056 30000
rect 7224 29600 7280 30000
rect 7448 29600 7504 30000
rect 7672 29600 7728 30000
rect 7896 29600 7952 30000
rect 8120 29600 8176 30000
rect 8344 29600 8400 30000
rect 8568 29600 8624 30000
rect 8792 29600 8848 30000
rect 9016 29600 9072 30000
rect 9240 29600 9296 30000
rect 9464 29600 9520 30000
rect 9688 29600 9744 30000
rect 9912 29600 9968 30000
rect 10136 29600 10192 30000
rect 10360 29600 10416 30000
rect 10584 29600 10640 30000
rect 10808 29600 10864 30000
rect 11032 29600 11088 30000
rect 11256 29600 11312 30000
rect 11480 29600 11536 30000
rect 11704 29600 11760 30000
rect 11928 29600 11984 30000
rect 12152 29600 12208 30000
rect 12376 29600 12432 30000
rect 12600 29600 12656 30000
rect 12824 29600 12880 30000
rect 13048 29600 13104 30000
rect 13272 29600 13328 30000
rect 13496 29600 13552 30000
rect 13720 29600 13776 30000
rect 13944 29600 14000 30000
rect 14168 29600 14224 30000
rect 14392 29600 14448 30000
rect 14616 29600 14672 30000
rect 14840 29600 14896 30000
rect 15064 29600 15120 30000
rect 15288 29600 15344 30000
rect 15512 29600 15568 30000
rect 15736 29600 15792 30000
rect 15960 29600 16016 30000
rect 16184 29600 16240 30000
rect 16408 29600 16464 30000
rect 16632 29600 16688 30000
rect 16856 29600 16912 30000
rect 17080 29600 17136 30000
rect 17304 29600 17360 30000
rect 17528 29600 17584 30000
rect 17752 29600 17808 30000
rect 17976 29600 18032 30000
rect 18200 29600 18256 30000
rect 18424 29600 18480 30000
rect 18648 29600 18704 30000
rect 18872 29600 18928 30000
rect 19096 29600 19152 30000
rect 19320 29600 19376 30000
rect 19544 29600 19600 30000
rect 19768 29600 19824 30000
rect 19992 29600 20048 30000
rect 20216 29600 20272 30000
rect 20440 29600 20496 30000
rect 20664 29600 20720 30000
rect 20888 29600 20944 30000
rect 21112 29600 21168 30000
rect 21336 29600 21392 30000
rect 21560 29600 21616 30000
rect 21784 29600 21840 30000
rect 22008 29600 22064 30000
rect 22232 29600 22288 30000
rect 22456 29600 22512 30000
rect 22680 29600 22736 30000
rect 22904 29600 22960 30000
rect 23128 29600 23184 30000
rect 23352 29600 23408 30000
rect 23576 29600 23632 30000
rect 23800 29600 23856 30000
rect 24024 29600 24080 30000
rect 24248 29600 24304 30000
rect 24472 29600 24528 30000
rect 24696 29600 24752 30000
rect 24920 29600 24976 30000
rect 25144 29600 25200 30000
rect 25368 29600 25424 30000
rect 25592 29600 25648 30000
rect 25816 29600 25872 30000
rect 26040 29600 26096 30000
rect 26264 29600 26320 30000
rect 26488 29600 26544 30000
rect 26712 29600 26768 30000
rect 26936 29600 26992 30000
rect 27160 29600 27216 30000
rect 27384 29600 27440 30000
rect 27608 29600 27664 30000
rect 7448 0 7504 400
rect 22400 0 22456 400
<< obsm2 >>
rect 2238 29570 2266 29600
rect 2382 29570 2490 29600
rect 2606 29570 2714 29600
rect 2830 29570 2938 29600
rect 3054 29570 3162 29600
rect 3278 29570 3386 29600
rect 3502 29570 3610 29600
rect 3726 29570 3834 29600
rect 3950 29570 4058 29600
rect 4174 29570 4282 29600
rect 4398 29570 4506 29600
rect 4622 29570 4730 29600
rect 4846 29570 4954 29600
rect 5070 29570 5178 29600
rect 5294 29570 5402 29600
rect 5518 29570 5626 29600
rect 5742 29570 5850 29600
rect 5966 29570 6074 29600
rect 6190 29570 6298 29600
rect 6414 29570 6522 29600
rect 6638 29570 6746 29600
rect 6862 29570 6970 29600
rect 7086 29570 7194 29600
rect 7310 29570 7418 29600
rect 7534 29570 7642 29600
rect 7758 29570 7866 29600
rect 7982 29570 8090 29600
rect 8206 29570 8314 29600
rect 8430 29570 8538 29600
rect 8654 29570 8762 29600
rect 8878 29570 8986 29600
rect 9102 29570 9210 29600
rect 9326 29570 9434 29600
rect 9550 29570 9658 29600
rect 9774 29570 9882 29600
rect 9998 29570 10106 29600
rect 10222 29570 10330 29600
rect 10446 29570 10554 29600
rect 10670 29570 10778 29600
rect 10894 29570 11002 29600
rect 11118 29570 11226 29600
rect 11342 29570 11450 29600
rect 11566 29570 11674 29600
rect 11790 29570 11898 29600
rect 12014 29570 12122 29600
rect 12238 29570 12346 29600
rect 12462 29570 12570 29600
rect 12686 29570 12794 29600
rect 12910 29570 13018 29600
rect 13134 29570 13242 29600
rect 13358 29570 13466 29600
rect 13582 29570 13690 29600
rect 13806 29570 13914 29600
rect 14030 29570 14138 29600
rect 14254 29570 14362 29600
rect 14478 29570 14586 29600
rect 14702 29570 14810 29600
rect 14926 29570 15034 29600
rect 15150 29570 15258 29600
rect 15374 29570 15482 29600
rect 15598 29570 15706 29600
rect 15822 29570 15930 29600
rect 16046 29570 16154 29600
rect 16270 29570 16378 29600
rect 16494 29570 16602 29600
rect 16718 29570 16826 29600
rect 16942 29570 17050 29600
rect 17166 29570 17274 29600
rect 17390 29570 17498 29600
rect 17614 29570 17722 29600
rect 17838 29570 17946 29600
rect 18062 29570 18170 29600
rect 18286 29570 18394 29600
rect 18510 29570 18618 29600
rect 18734 29570 18842 29600
rect 18958 29570 19066 29600
rect 19182 29570 19290 29600
rect 19406 29570 19514 29600
rect 19630 29570 19738 29600
rect 19854 29570 19962 29600
rect 20078 29570 20186 29600
rect 20302 29570 20410 29600
rect 20526 29570 20634 29600
rect 20750 29570 20858 29600
rect 20974 29570 21082 29600
rect 21198 29570 21306 29600
rect 21422 29570 21530 29600
rect 21646 29570 21754 29600
rect 21870 29570 21978 29600
rect 22094 29570 22202 29600
rect 22318 29570 22426 29600
rect 22542 29570 22650 29600
rect 22766 29570 22874 29600
rect 22990 29570 23098 29600
rect 23214 29570 23322 29600
rect 23438 29570 23546 29600
rect 23662 29570 23770 29600
rect 23886 29570 23994 29600
rect 24110 29570 24218 29600
rect 24334 29570 24442 29600
rect 24558 29570 24666 29600
rect 24782 29570 24890 29600
rect 25006 29570 25114 29600
rect 25230 29570 25338 29600
rect 25454 29570 25562 29600
rect 25678 29570 25786 29600
rect 25902 29570 26010 29600
rect 26126 29570 26234 29600
rect 26350 29570 26458 29600
rect 26574 29570 26682 29600
rect 26798 29570 26906 29600
rect 27022 29570 27130 29600
rect 27246 29570 27354 29600
rect 27470 29570 27578 29600
rect 27694 29570 27762 29600
rect 2238 1549 27762 29570
<< obsm3 >>
rect 2233 1554 27767 28322
<< metal4 >>
rect 2224 1538 2384 28254
rect 9904 1538 10064 28254
rect 17584 1538 17744 28254
rect 25264 1538 25424 28254
<< labels >>
rlabel metal2 s 2296 29600 2352 30000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 9016 29600 9072 30000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 9688 29600 9744 30000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 10360 29600 10416 30000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 11032 29600 11088 30000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 11704 29600 11760 30000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 12376 29600 12432 30000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 13048 29600 13104 30000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 13720 29600 13776 30000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 14392 29600 14448 30000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 15064 29600 15120 30000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 2968 29600 3024 30000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 15736 29600 15792 30000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 16408 29600 16464 30000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 17080 29600 17136 30000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 17752 29600 17808 30000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 18424 29600 18480 30000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 19096 29600 19152 30000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 19768 29600 19824 30000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 20440 29600 20496 30000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 21112 29600 21168 30000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 21784 29600 21840 30000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 3640 29600 3696 30000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 22456 29600 22512 30000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 23128 29600 23184 30000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 23800 29600 23856 30000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 24472 29600 24528 30000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 25144 29600 25200 30000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 25816 29600 25872 30000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 26488 29600 26544 30000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 27160 29600 27216 30000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 4312 29600 4368 30000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 4984 29600 5040 30000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 5656 29600 5712 30000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 6328 29600 6384 30000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 7000 29600 7056 30000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 7672 29600 7728 30000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 8344 29600 8400 30000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2520 29600 2576 30000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 9240 29600 9296 30000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 9912 29600 9968 30000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 10584 29600 10640 30000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 11256 29600 11312 30000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 11928 29600 11984 30000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 12600 29600 12656 30000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 13272 29600 13328 30000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 13944 29600 14000 30000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 14616 29600 14672 30000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 15288 29600 15344 30000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3192 29600 3248 30000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 15960 29600 16016 30000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 16632 29600 16688 30000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 17304 29600 17360 30000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 17976 29600 18032 30000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 18648 29600 18704 30000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 19320 29600 19376 30000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 19992 29600 20048 30000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 20664 29600 20720 30000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 21336 29600 21392 30000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 22008 29600 22064 30000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 3864 29600 3920 30000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 22680 29600 22736 30000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 23352 29600 23408 30000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 24024 29600 24080 30000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 24696 29600 24752 30000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 25368 29600 25424 30000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 26040 29600 26096 30000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 26712 29600 26768 30000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 27384 29600 27440 30000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 4536 29600 4592 30000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 5208 29600 5264 30000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 5880 29600 5936 30000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 6552 29600 6608 30000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 7224 29600 7280 30000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 7896 29600 7952 30000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 8568 29600 8624 30000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2744 29600 2800 30000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 9464 29600 9520 30000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 10136 29600 10192 30000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 10808 29600 10864 30000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 11480 29600 11536 30000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 12152 29600 12208 30000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 12824 29600 12880 30000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 13496 29600 13552 30000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 14168 29600 14224 30000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 14840 29600 14896 30000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 15512 29600 15568 30000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 3416 29600 3472 30000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 16184 29600 16240 30000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 16856 29600 16912 30000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 17528 29600 17584 30000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 18200 29600 18256 30000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 18872 29600 18928 30000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 19544 29600 19600 30000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 20216 29600 20272 30000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 20888 29600 20944 30000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 21560 29600 21616 30000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 22232 29600 22288 30000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 4088 29600 4144 30000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 22904 29600 22960 30000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 23576 29600 23632 30000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 24248 29600 24304 30000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 24920 29600 24976 30000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 25592 29600 25648 30000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 26264 29600 26320 30000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 26936 29600 26992 30000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 27608 29600 27664 30000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 4760 29600 4816 30000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 5432 29600 5488 30000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 6104 29600 6160 30000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 6776 29600 6832 30000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 7448 29600 7504 30000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 8120 29600 8176 30000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 8792 29600 8848 30000 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 2224 1538 2384 28254 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 28254 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 28254 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 28254 6 vss
port 116 nsew ground bidirectional
rlabel metal2 s 7448 0 7504 400 6 wb_clk_i
port 117 nsew signal input
rlabel metal2 s 22400 0 22456 400 6 wb_rst_i
port 118 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 420296
string GDS_FILE /home/mm4uz/asic/gf180-shuttle-0/submission/gf180-ceylanM/openlane/wrapped_multiplier_8/runs/22_12_05_17_33/results/signoff/wrapped_multiplier_8.magic.gds
string GDS_START 50130
<< end >>

